// -----------------------------------------------------------------------------
//
// -----------------------------------------------------------------------------
// Description:
// ------------
//
// CSD borrow save representation to two's complement conversion.
//
// -----------------------------------------------------------------------------
// File name:
// ----------
//
// csd2bin.v
//
// -----------------------------------------------------------------------------
// Interface:
// ----------
//
//  Clock, reset & enable inputs:
//    - None
//
//  Data inputs:
//    - x         : X input variable (two's complement, W bits).
//
//  Data outputs:
//    - y         : Y output result (cannonic signed digit, 2*W bits).
//
//  Parameters:
//    - W         : Word width (natural, default: 64).
//
// -----------------------------------------------------------------------------
// History:
// --------
//
//    - 2016-04-18 - ilesser - Original version.
//
// -----------------------------------------------------------------------------

// *****************************************************************************
// Interface
// *****************************************************************************
module csd2bin #(
    // ----------------------------------
    // Parameters
    // ----------------------------------
    parameter W      = 64
  ) (
    // ----------------------------------
    // Data inputs
    // ----------------------------------
    input   wire  [2*W-1:0]   x,
    // ----------------------------------
    // Data outputs
    // ----------------------------------
    output  reg   [W-1:0]     y
  );
// *****************************************************************************

// *****************************************************************************
// Architecture
// *****************************************************************************
//    x_i = {x_i^s x_i^d}
//
//    y_i = x_i^d - x_i^s
//
//    y   = x^d - x^s = x^d + ~x^s + '1'
//
// *****************************************************************************
//
//
//                x
//                 i
//                | |
//                O |
//              +-----+
//              |     |
//     c -------| FA  |------ c        c  = 1'b1
//      i+1     |     |        i        0
//              +-----+
//                 |
//                 |
//                 |
//                 |
//                 y
//                  i
//
//
//       +-----------+----------+
//       |    ci=0   |    ci=1  |
//  +----+------+----+------+---+
//  | xi | ci+1 |si  | ci+1 |si |
//  +----+------+----+------+---+
//  | 00 |  0   | 1  |  1   | 0 |
//  | 01 |  1   | 0  |  1   | 1 |
//  | 10 |  0   | 0  |  0   | 1 |
//  | 11 |  0   | 1  |  1   | 0 |
//  +----+------+----+------+---+
//
// *****************************************************************************


   // -----------------------------------------------------
   // Internal signals
   // -----------------------------------------------------
   reg   [W:0]       c;    // carry
   reg   [W-1:0]     x_s;  // x sign bit
   reg   [W-1:0]     x_d;  // x data bit
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Combinational logic
   // -----------------------------------------------------
   //always @(*) begin
   //   c[0] = 1'b1;
   //end
   assign c[0] = 1'b1;

   genvar i;
   generate
      for (i=0; i < W; i=i+1) begin
         always @(*) begin

            // Split the CSD numbers into its BS representation
            // _s stands for sign bit and _d for data bit
            {x_s[i], x_d[i]}  = x[2*i+1:2*i];

            // Propagate the carry
            {c[i+1], y[i]}    = !x_s[i] + x_d[i] + c[i];

         end
      end
   endgenerate
   // -----------------------------------------------------

// *****************************************************************************

// *****************************************************************************
// Assertions and debugging
// *****************************************************************************
`ifdef RTL_DEBUG

   //XXXXX TO FILL IN HERE XXXXX

`endif
// *****************************************************************************

endmodule

