//--------------------------------------------------------------------------------
//
// BKM LUT automatically generated on 06:12:19 PM (ART) Wednesday 31 August 2016
// using the bkm_lut.m function. Version = 1.0, from Monday 29 August 2016.
// Parameters:
// Number of steps of the algorithm:   N  = 64
// Word size of the data channel:      WD = 73
// Word size of the control channel:   WC = 21
// Integer word size:                  WI = 11
//
//--------------------------------------------------------------------------------
assign X[4'b0000] [00] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-1+1) + ( 0^2+ 0^2) * 2^(-2*1) )   n =  1   d_n = 0 
assign X[4'b0000] [01] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-2+1) + ( 0^2+ 0^2) * 2^(-2*2) )   n =  2   d_n = 0 
assign X[4'b0000] [02] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-3+1) + ( 0^2+ 0^2) * 2^(-2*3) )   n =  3   d_n = 0 
assign X[4'b0000] [03] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-4+1) + ( 0^2+ 0^2) * 2^(-2*4) )   n =  4   d_n = 0 
assign X[4'b0000] [04] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-5+1) + ( 0^2+ 0^2) * 2^(-2*5) )   n =  5   d_n = 0 
assign X[4'b0000] [05] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-6+1) + ( 0^2+ 0^2) * 2^(-2*6) )   n =  6   d_n = 0 
assign X[4'b0000] [06] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-7+1) + ( 0^2+ 0^2) * 2^(-2*7) )   n =  7   d_n = 0 
assign X[4'b0000] [07] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-8+1) + ( 0^2+ 0^2) * 2^(-2*8) )   n =  8   d_n = 0 
assign X[4'b0000] [08] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-9+1) + ( 0^2+ 0^2) * 2^(-2*9) )   n =  9   d_n = 0 
assign X[4'b0000] [09] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = 0 
assign X[4'b0000] [10] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = 0 
assign X[4'b0000] [11] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = 0 
assign X[4'b0000] [12] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = 0 
assign X[4'b0000] [13] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = 0 
assign X[4'b0000] [14] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = 0 
assign X[4'b0000] [15] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = 0 
assign X[4'b0000] [16] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = 0 
assign X[4'b0000] [17] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = 0 
assign X[4'b0000] [18] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = 0 
assign X[4'b0000] [19] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = 0 
assign X[4'b0000] [20] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = 0 
assign X[4'b0000] [21] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = 0 
assign X[4'b0000] [22] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = 0 
assign X[4'b0000] [23] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = 0 
assign X[4'b0000] [24] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = 0 
assign X[4'b0000] [25] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = 0 
assign X[4'b0000] [26] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = 0 
assign X[4'b0000] [27] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = 0 
assign X[4'b0000] [28] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = 0 
assign X[4'b0000] [29] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = 0 
assign X[4'b0000] [30] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = 0 
assign X[4'b0000] [31] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = 0 
assign X[4'b0000] [32] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = 0 
assign X[4'b0000] [33] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = 0 
assign X[4'b0000] [34] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = 0 
assign X[4'b0000] [35] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = 0 
assign X[4'b0000] [36] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = 0 
assign X[4'b0000] [37] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = 0 
assign X[4'b0000] [38] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = 0 
assign X[4'b0000] [39] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = 0 
assign X[4'b0000] [40] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = 0 
assign X[4'b0000] [41] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = 0 
assign X[4'b0000] [42] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = 0 
assign X[4'b0000] [43] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = 0 
assign X[4'b0000] [44] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = 0 
assign X[4'b0000] [45] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = 0 
assign X[4'b0000] [46] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = 0 
assign X[4'b0000] [47] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = 0 
assign X[4'b0000] [48] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = 0 
assign X[4'b0000] [49] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = 0 
assign X[4'b0000] [50] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = 0 
assign X[4'b0000] [51] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = 0 
assign X[4'b0000] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = 0 
assign X[4'b0000] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = 0 
assign X[4'b0000] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = 0 
assign X[4'b0000] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = 0 
assign X[4'b0000] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = 0 
assign X[4'b0000] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = 0 
assign X[4'b0000] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = 0 
assign X[4'b0000] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = 0 
assign X[4'b0000] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = 0 
assign X[4'b0000] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = 0 
assign X[4'b0000] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = 0 
assign X[4'b0000] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = 0 
assign X[4'b0001] [00] = 146'h 0000004C40313041003400000000000000000;  // +0.4054651081081644 = 0.5 * ln( 1 +  1 * 2^(-1+1) + ( 1^2+ 0^2) * 2^(-2*1) )   n =  1   d_n = 1 
assign X[4'b0001] [01] = 146'h 00000010C104000300C100000000000000000;  // +0.2231435513142098 = 0.5 * ln( 1 +  1 * 2^(-2+1) + ( 1^2+ 0^2) * 2^(-2*2) )   n =  2   d_n = 1 
assign X[4'b0001] [02] = 146'h 000000040C04430040C300000000000000000;  // +0.1177830356563835 = 0.5 * ln( 1 +  1 * 2^(-3+1) + ( 1^2+ 0^2) * 2^(-2*3) )   n =  3   d_n = 1 
assign X[4'b0001] [03] = 146'h 0000000100C01104C04C00000000000000000;  // +0.0606246218164348 = 0.5 * ln( 1 +  1 * 2^(-4+1) + ( 1^2+ 0^2) * 2^(-2*4) )   n =  4   d_n = 1 
assign X[4'b0001] [04] = 146'h 00000000400C0044433010000000000000000;  // +0.0307716586667537 = 0.5 * ln( 1 +  1 * 2^(-5+1) + ( 1^2+ 0^2) * 2^(-2*5) )   n =  5   d_n = 1 
assign X[4'b0001] [05] = 146'h 000000001000C0011104CC000000000000000;  // +0.0155041865359653 = 0.5 * ln( 1 +  1 * 2^(-6+1) + ( 1^2+ 0^2) * 2^(-2*6) )   n =  6   d_n = 1 
assign X[4'b0001] [06] = 146'h 0000000004000C00044443400000000000000;  // +0.0077821404420549 = 0.5 * ln( 1 +  1 * 2^(-7+1) + ( 1^2+ 0^2) * 2^(-2*7) )   n =  7   d_n = 1 
assign X[4'b0001] [07] = 146'h 00000000010000C0001111000000000000000;  // +0.0038986404156573 = 0.5 * ln( 1 +  1 * 2^(-8+1) + ( 1^2+ 0^2) * 2^(-2*8) )   n =  8   d_n = 1 
assign X[4'b0001] [08] = 146'h 000000000040000C000044440000000000000;  // +0.0019512201312617 = 0.5 * ln( 1 +  1 * 2^(-9+1) + ( 1^2+ 0^2) * 2^(-2*9) )   n =  9   d_n = 1 
assign X[4'b0001] [09] = 146'h 0000000000100000C00001110000000000000;  // +0.0009760859730555 = 0.5 * ln( 1 +  1 * 2^(-10+1) + ( 1^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = 1 
assign X[4'b0001] [10] = 146'h 00000000000400000C0000044000000000000;  // +0.0004881620795014 = 0.5 * ln( 1 +  1 * 2^(-11+1) + ( 1^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = 1 
assign X[4'b0001] [11] = 146'h 000000000001000000C000001000000000000;  // +0.0002441108275274 = 0.5 * ln( 1 +  1 * 2^(-12+1) + ( 1^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = 1 
assign X[4'b0001] [12] = 146'h 0000000000004000000C00000000000000000;  // +0.0001220628625257 = 0.5 * ln( 1 +  1 * 2^(-13+1) + ( 1^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = 1 
assign X[4'b0001] [13] = 146'h 00000000000010000000C0000000000000000;  // +0.0000610332936806 = 0.5 * ln( 1 +  1 * 2^(-14+1) + ( 1^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = 1 
assign X[4'b0001] [14] = 146'h 000000000000040000000C000000000000000;  // +0.0000305171124732 = 0.5 * ln( 1 +  1 * 2^(-15+1) + ( 1^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = 1 
assign X[4'b0001] [15] = 146'h 0000000000000100000000C00000000000000;  // +0.0000152586726484 = 0.5 * ln( 1 +  1 * 2^(-16+1) + ( 1^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = 1 
assign X[4'b0001] [16] = 146'h 00000000000000400000000C0000000000000;  // +0.0000076293654276 = 0.5 * ln( 1 +  1 * 2^(-17+1) + ( 1^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = 1 
assign X[4'b0001] [17] = 146'h 000000000000001000000000C000000000000;  // +0.0000038146899897 = 0.5 * ln( 1 +  1 * 2^(-18+1) + ( 1^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = 1 
assign X[4'b0001] [18] = 146'h 0000000000000004000000000C00000000000;  // +0.0000019073468138 = 0.5 * ln( 1 +  1 * 2^(-19+1) + ( 1^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = 1 
assign X[4'b0001] [19] = 146'h 00000000000000010000000000C0000000000;  // +0.0000009536738617 = 0.5 * ln( 1 +  1 * 2^(-20+1) + ( 1^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = 1 
assign X[4'b0001] [20] = 146'h 000000000000000040000000000C000000000;  // +0.0000004768370445 = 0.5 * ln( 1 +  1 * 2^(-21+1) + ( 1^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = 1 
assign X[4'b0001] [21] = 146'h 0000000000000000100000000000C00000000;  // +0.0000002384185507 = 0.5 * ln( 1 +  1 * 2^(-22+1) + ( 1^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = 1 
assign X[4'b0001] [22] = 146'h 00000000000000000400000000000C0000000;  // +0.0000001192092824 = 0.5 * ln( 1 +  1 * 2^(-23+1) + ( 1^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = 1 
assign X[4'b0001] [23] = 146'h 000000000000000001000000000000C000000;  // +0.0000000596046430 = 0.5 * ln( 1 +  1 * 2^(-24+1) + ( 1^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = 1 
assign X[4'b0001] [24] = 146'h 0000000000000000004000000000000C00000;  // +0.0000000298023219 = 0.5 * ln( 1 +  1 * 2^(-25+1) + ( 1^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = 1 
assign X[4'b0001] [25] = 146'h 0000000000000000001000000000000100000;  // +0.0000000149011611 = 0.5 * ln( 1 +  1 * 2^(-26+1) + ( 1^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = 1 
assign X[4'b0001] [26] = 146'h 0000000000000000000400000000000000000;  // +0.0000000074505806 = 0.5 * ln( 1 +  1 * 2^(-27+1) + ( 1^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = 1 
assign X[4'b0001] [27] = 146'h 0000000000000000000100000000000000000;  // +0.0000000037252903 = 0.5 * ln( 1 +  1 * 2^(-28+1) + ( 1^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = 1 
assign X[4'b0001] [28] = 146'h 0000000000000000000040000000000000000;  // +0.0000000018626451 = 0.5 * ln( 1 +  1 * 2^(-29+1) + ( 1^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = 1 
assign X[4'b0001] [29] = 146'h 0000000000000000000010000000000000000;  // +0.0000000009313226 = 0.5 * ln( 1 +  1 * 2^(-30+1) + ( 1^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = 1 
assign X[4'b0001] [30] = 146'h 0000000000000000000004000000000000000;  // +0.0000000004656613 = 0.5 * ln( 1 +  1 * 2^(-31+1) + ( 1^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = 1 
assign X[4'b0001] [31] = 146'h 0000000000000000000001000000000000000;  // +0.0000000002328306 = 0.5 * ln( 1 +  1 * 2^(-32+1) + ( 1^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = 1 
assign X[4'b0001] [32] = 146'h 0000000000000000000000400000000000000;  // +0.0000000001164153 = 0.5 * ln( 1 +  1 * 2^(-33+1) + ( 1^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = 1 
assign X[4'b0001] [33] = 146'h 0000000000000000000000100000000000000;  // +0.0000000000582077 = 0.5 * ln( 1 +  1 * 2^(-34+1) + ( 1^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = 1 
assign X[4'b0001] [34] = 146'h 0000000000000000000000040000000000000;  // +0.0000000000291038 = 0.5 * ln( 1 +  1 * 2^(-35+1) + ( 1^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = 1 
assign X[4'b0001] [35] = 146'h 0000000000000000000000010000000000000;  // +0.0000000000145519 = 0.5 * ln( 1 +  1 * 2^(-36+1) + ( 1^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = 1 
assign X[4'b0001] [36] = 146'h 0000000000000000000000004000000000000;  // +0.0000000000072760 = 0.5 * ln( 1 +  1 * 2^(-37+1) + ( 1^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = 1 
assign X[4'b0001] [37] = 146'h 0000000000000000000000001000000000000;  // +0.0000000000036380 = 0.5 * ln( 1 +  1 * 2^(-38+1) + ( 1^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = 1 
assign X[4'b0001] [38] = 146'h 0000000000000000000000000400000000000;  // +0.0000000000018190 = 0.5 * ln( 1 +  1 * 2^(-39+1) + ( 1^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = 1 
assign X[4'b0001] [39] = 146'h 0000000000000000000000000100000000000;  // +0.0000000000009095 = 0.5 * ln( 1 +  1 * 2^(-40+1) + ( 1^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = 1 
assign X[4'b0001] [40] = 146'h 0000000000000000000000000040000000000;  // +0.0000000000004547 = 0.5 * ln( 1 +  1 * 2^(-41+1) + ( 1^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = 1 
assign X[4'b0001] [41] = 146'h 0000000000000000000000000010000000000;  // +0.0000000000002274 = 0.5 * ln( 1 +  1 * 2^(-42+1) + ( 1^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = 1 
assign X[4'b0001] [42] = 146'h 0000000000000000000000000004000000000;  // +0.0000000000001137 = 0.5 * ln( 1 +  1 * 2^(-43+1) + ( 1^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = 1 
assign X[4'b0001] [43] = 146'h 0000000000000000000000000001000000000;  // +0.0000000000000568 = 0.5 * ln( 1 +  1 * 2^(-44+1) + ( 1^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = 1 
assign X[4'b0001] [44] = 146'h 0000000000000000000000000000400000000;  // +0.0000000000000284 = 0.5 * ln( 1 +  1 * 2^(-45+1) + ( 1^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = 1 
assign X[4'b0001] [45] = 146'h 0000000000000000000000000000100000000;  // +0.0000000000000142 = 0.5 * ln( 1 +  1 * 2^(-46+1) + ( 1^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = 1 
assign X[4'b0001] [46] = 146'h 0000000000000000000000000000040000000;  // +0.0000000000000071 = 0.5 * ln( 1 +  1 * 2^(-47+1) + ( 1^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = 1 
assign X[4'b0001] [47] = 146'h 0000000000000000000000000000010000000;  // +0.0000000000000036 = 0.5 * ln( 1 +  1 * 2^(-48+1) + ( 1^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = 1 
assign X[4'b0001] [48] = 146'h 0000000000000000000000000000004000000;  // +0.0000000000000018 = 0.5 * ln( 1 +  1 * 2^(-49+1) + ( 1^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = 1 
assign X[4'b0001] [49] = 146'h 0000000000000000000000000000001000000;  // +0.0000000000000009 = 0.5 * ln( 1 +  1 * 2^(-50+1) + ( 1^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = 1 
assign X[4'b0001] [50] = 146'h 0000000000000000000000000000000400000;  // +0.0000000000000004 = 0.5 * ln( 1 +  1 * 2^(-51+1) + ( 1^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = 1 
assign X[4'b0001] [51] = 146'h 0000000000000000000000000000000100000;  // +0.0000000000000002 = 0.5 * ln( 1 +  1 * 2^(-52+1) + ( 1^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = 1 
assign X[4'b0001] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-53+1) + ( 1^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = 1 
assign X[4'b0001] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-54+1) + ( 1^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = 1 
assign X[4'b0001] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-55+1) + ( 1^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = 1 
assign X[4'b0001] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-56+1) + ( 1^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = 1 
assign X[4'b0001] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-57+1) + ( 1^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = 1 
assign X[4'b0001] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-58+1) + ( 1^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = 1 
assign X[4'b0001] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-59+1) + ( 1^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = 1 
assign X[4'b0001] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-60+1) + ( 1^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = 1 
assign X[4'b0001] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-61+1) + ( 1^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = 1 
assign X[4'b0001] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-62+1) + ( 1^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = 1 
assign X[4'b0001] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-63+1) + ( 1^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = 1 
assign X[4'b0001] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-64+1) + ( 1^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = 1 
assign X[4'b0010] [00] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-1+1) + ( 0^2+ 0^2) * 2^(-2*1) )   n =  1   d_n = -0 
assign X[4'b0010] [01] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-2+1) + ( 0^2+ 0^2) * 2^(-2*2) )   n =  2   d_n = -0 
assign X[4'b0010] [02] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-3+1) + ( 0^2+ 0^2) * 2^(-2*3) )   n =  3   d_n = -0 
assign X[4'b0010] [03] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-4+1) + ( 0^2+ 0^2) * 2^(-2*4) )   n =  4   d_n = -0 
assign X[4'b0010] [04] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-5+1) + ( 0^2+ 0^2) * 2^(-2*5) )   n =  5   d_n = -0 
assign X[4'b0010] [05] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-6+1) + ( 0^2+ 0^2) * 2^(-2*6) )   n =  6   d_n = -0 
assign X[4'b0010] [06] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-7+1) + ( 0^2+ 0^2) * 2^(-2*7) )   n =  7   d_n = -0 
assign X[4'b0010] [07] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-8+1) + ( 0^2+ 0^2) * 2^(-2*8) )   n =  8   d_n = -0 
assign X[4'b0010] [08] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-9+1) + ( 0^2+ 0^2) * 2^(-2*9) )   n =  9   d_n = -0 
assign X[4'b0010] [09] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = -0 
assign X[4'b0010] [10] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = -0 
assign X[4'b0010] [11] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = -0 
assign X[4'b0010] [12] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = -0 
assign X[4'b0010] [13] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = -0 
assign X[4'b0010] [14] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = -0 
assign X[4'b0010] [15] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = -0 
assign X[4'b0010] [16] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = -0 
assign X[4'b0010] [17] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = -0 
assign X[4'b0010] [18] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = -0 
assign X[4'b0010] [19] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = -0 
assign X[4'b0010] [20] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = -0 
assign X[4'b0010] [21] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = -0 
assign X[4'b0010] [22] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = -0 
assign X[4'b0010] [23] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = -0 
assign X[4'b0010] [24] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = -0 
assign X[4'b0010] [25] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = -0 
assign X[4'b0010] [26] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = -0 
assign X[4'b0010] [27] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = -0 
assign X[4'b0010] [28] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = -0 
assign X[4'b0010] [29] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = -0 
assign X[4'b0010] [30] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = -0 
assign X[4'b0010] [31] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = -0 
assign X[4'b0010] [32] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = -0 
assign X[4'b0010] [33] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = -0 
assign X[4'b0010] [34] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = -0 
assign X[4'b0010] [35] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = -0 
assign X[4'b0010] [36] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = -0 
assign X[4'b0010] [37] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = -0 
assign X[4'b0010] [38] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = -0 
assign X[4'b0010] [39] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = -0 
assign X[4'b0010] [40] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = -0 
assign X[4'b0010] [41] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = -0 
assign X[4'b0010] [42] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = -0 
assign X[4'b0010] [43] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = -0 
assign X[4'b0010] [44] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = -0 
assign X[4'b0010] [45] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = -0 
assign X[4'b0010] [46] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = -0 
assign X[4'b0010] [47] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = -0 
assign X[4'b0010] [48] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = -0 
assign X[4'b0010] [49] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = -0 
assign X[4'b0010] [50] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = -0 
assign X[4'b0010] [51] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = -0 
assign X[4'b0010] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = -0 
assign X[4'b0010] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = -0 
assign X[4'b0010] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = -0 
assign X[4'b0010] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = -0 
assign X[4'b0010] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = -0 
assign X[4'b0010] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = -0 
assign X[4'b0010] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = -0 
assign X[4'b0010] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = -0 
assign X[4'b0010] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = -0 
assign X[4'b0010] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = -0 
assign X[4'b0010] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = -0 
assign X[4'b0010] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = -0 
assign X[4'b0011] [00] = 146'h 000003110C410C0C400000000000000000000;  // -0.6931471805599453 = 0.5 * ln( 1 + -1 * 2^(-1+1) + (-1^2+ 0^2) * 2^(-2*1) )   n =  1   d_n = -1 
assign X[4'b0011] [01] = 146'h 00000030CC4CC440C03000000000000000000;  // -0.2876820724517809 = 0.5 * ln( 1 + -1 * 2^(-2+1) + (-1^2+ 0^2) * 2^(-2*2) )   n =  2   d_n = -1 
assign X[4'b0011] [02] = 146'h 0000000C0C31010C130000000000000000000;  // -0.1335313926245226 = 0.5 * ln( 1 + -1 * 2^(-3+1) + (-1^2+ 0^2) * 2^(-2*3) )   n =  3   d_n = -1 
assign X[4'b0011] [03] = 146'h 0000000300C0C44C431040000000000000000;  // -0.0645385211375712 = 0.5 * ln( 1 + -1 * 2^(-4+1) + (-1^2+ 0^2) * 2^(-2*4) )   n =  4   d_n = -1 
assign X[4'b0011] [04] = 146'h 00000000C00C0311011030000000000000000;  // -0.0317486983145803 = 0.5 * ln( 1 + -1 * 2^(-5+1) + (-1^2+ 0^2) * 2^(-2*5) )   n =  5   d_n = -1 
assign X[4'b0011] [05] = 146'h 000000003000C00C444C44000000000000000;  // -0.0157483569681392 = 0.5 * ln( 1 + -1 * 2^(-6+1) + (-1^2+ 0^2) * 2^(-2*6) )   n =  6   d_n = -1 
assign X[4'b0011] [06] = 146'h 000000000C000C00311101000000000000000;  // -0.0078431774610259 = 0.5 * ln( 1 + -1 * 2^(-7+1) + (-1^2+ 0^2) * 2^(-2*7) )   n =  7   d_n = -1 
assign X[4'b0011] [07] = 146'h 00000000030000C000C444400000000000000;  // -0.0039138993211363 = 0.5 * ln( 1 + -1 * 2^(-8+1) + (-1^2+ 0^2) * 2^(-2*8) )   n =  8   d_n = -1 
assign X[4'b0011] [08] = 146'h 0000000000C0000C000311100000000000000;  // -0.0019550348358034 = 0.5 * ln( 1 + -1 * 2^(-9+1) + (-1^2+ 0^2) * 2^(-2*9) )   n =  9   d_n = -1 
assign X[4'b0011] [09] = 146'h 0000000000300000C0000C440000000000000;  // -0.0009770396478266 = 0.5 * ln( 1 + -1 * 2^(-10+1) + (-1^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = -1 
assign X[4'b0011] [10] = 146'h 00000000000C00000C0000310000000000000;  // -0.0004884004981089 = 0.5 * ln( 1 + -1 * 2^(-11+1) + (-1^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = -1 
assign X[4'b0011] [11] = 146'h 000000000003000000C00000C000000000000;  // -0.0002441704321739 = 0.5 * ln( 1 + -1 * 2^(-12+1) + (-1^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = -1 
assign X[4'b0011] [12] = 146'h 000000000000C000000C00000000000000000;  // -0.0001220777636870 = 0.5 * ln( 1 + -1 * 2^(-13+1) + (-1^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = -1 
assign X[4'b0011] [13] = 146'h 00000000000030000000C0000000000000000;  // -0.0000610370189709 = 0.5 * ln( 1 + -1 * 2^(-14+1) + (-1^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = -1 
assign X[4'b0011] [14] = 146'h 0000000000000C0000000C000000000000000;  // -0.0000305180437958 = 0.5 * ln( 1 + -1 * 2^(-15+1) + (-1^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = -1 
assign X[4'b0011] [15] = 146'h 0000000000000300000000C00000000000000;  // -0.0000152589054790 = 0.5 * ln( 1 + -1 * 2^(-16+1) + (-1^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = -1 
assign X[4'b0011] [16] = 146'h 00000000000000C00000000C0000000000000;  // -0.0000076294236352 = 0.5 * ln( 1 + -1 * 2^(-17+1) + (-1^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = -1 
assign X[4'b0011] [17] = 146'h 000000000000003000000000C000000000000;  // -0.0000038147045416 = 0.5 * ln( 1 + -1 * 2^(-18+1) + (-1^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = -1 
assign X[4'b0011] [18] = 146'h 000000000000000C000000000C00000000000;  // -0.0000019073504518 = 0.5 * ln( 1 + -1 * 2^(-19+1) + (-1^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = -1 
assign X[4'b0011] [19] = 146'h 00000000000000030000000000C0000000000;  // -0.0000009536747712 = 0.5 * ln( 1 + -1 * 2^(-20+1) + (-1^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = -1 
assign X[4'b0011] [20] = 146'h 0000000000000000C0000000000C000000000;  // -0.0000004768372719 = 0.5 * ln( 1 + -1 * 2^(-21+1) + (-1^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = -1 
assign X[4'b0011] [21] = 146'h 0000000000000000300000000000C00000000;  // -0.0000002384186075 = 0.5 * ln( 1 + -1 * 2^(-22+1) + (-1^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = -1 
assign X[4'b0011] [22] = 146'h 00000000000000000C00000000000C0000000;  // -0.0000001192092967 = 0.5 * ln( 1 + -1 * 2^(-23+1) + (-1^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = -1 
assign X[4'b0011] [23] = 146'h 000000000000000003000000000000C000000;  // -0.0000000596046466 = 0.5 * ln( 1 + -1 * 2^(-24+1) + (-1^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = -1 
assign X[4'b0011] [24] = 146'h 000000000000000000C000000000001000000;  // -0.0000000298023228 = 0.5 * ln( 1 + -1 * 2^(-25+1) + (-1^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = -1 
assign X[4'b0011] [25] = 146'h 0000000000000000003000000000000000000;  // -0.0000000149011613 = 0.5 * ln( 1 + -1 * 2^(-26+1) + (-1^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = -1 
assign X[4'b0011] [26] = 146'h 0000000000000000000C00000000000000000;  // -0.0000000074505806 = 0.5 * ln( 1 + -1 * 2^(-27+1) + (-1^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = -1 
assign X[4'b0011] [27] = 146'h 0000000000000000000300000000000000000;  // -0.0000000037252903 = 0.5 * ln( 1 + -1 * 2^(-28+1) + (-1^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = -1 
assign X[4'b0011] [28] = 146'h 00000000000000000000C0000000000000000;  // -0.0000000018626452 = 0.5 * ln( 1 + -1 * 2^(-29+1) + (-1^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = -1 
assign X[4'b0011] [29] = 146'h 0000000000000000000030000000000000000;  // -0.0000000009313226 = 0.5 * ln( 1 + -1 * 2^(-30+1) + (-1^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = -1 
assign X[4'b0011] [30] = 146'h 000000000000000000000C000000000000000;  // -0.0000000004656613 = 0.5 * ln( 1 + -1 * 2^(-31+1) + (-1^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = -1 
assign X[4'b0011] [31] = 146'h 0000000000000000000003000000000000000;  // -0.0000000002328306 = 0.5 * ln( 1 + -1 * 2^(-32+1) + (-1^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = -1 
assign X[4'b0011] [32] = 146'h 0000000000000000000000C00000000000000;  // -0.0000000001164153 = 0.5 * ln( 1 + -1 * 2^(-33+1) + (-1^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = -1 
assign X[4'b0011] [33] = 146'h 0000000000000000000000300000000000000;  // -0.0000000000582077 = 0.5 * ln( 1 + -1 * 2^(-34+1) + (-1^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = -1 
assign X[4'b0011] [34] = 146'h 00000000000000000000000C0000000000000;  // -0.0000000000291038 = 0.5 * ln( 1 + -1 * 2^(-35+1) + (-1^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = -1 
assign X[4'b0011] [35] = 146'h 0000000000000000000000030000000000000;  // -0.0000000000145519 = 0.5 * ln( 1 + -1 * 2^(-36+1) + (-1^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = -1 
assign X[4'b0011] [36] = 146'h 000000000000000000000000C000000000000;  // -0.0000000000072760 = 0.5 * ln( 1 + -1 * 2^(-37+1) + (-1^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = -1 
assign X[4'b0011] [37] = 146'h 0000000000000000000000003000000000000;  // -0.0000000000036380 = 0.5 * ln( 1 + -1 * 2^(-38+1) + (-1^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = -1 
assign X[4'b0011] [38] = 146'h 0000000000000000000000000C00000000000;  // -0.0000000000018190 = 0.5 * ln( 1 + -1 * 2^(-39+1) + (-1^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = -1 
assign X[4'b0011] [39] = 146'h 0000000000000000000000000300000000000;  // -0.0000000000009095 = 0.5 * ln( 1 + -1 * 2^(-40+1) + (-1^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = -1 
assign X[4'b0011] [40] = 146'h 00000000000000000000000000C0000000000;  // -0.0000000000004547 = 0.5 * ln( 1 + -1 * 2^(-41+1) + (-1^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = -1 
assign X[4'b0011] [41] = 146'h 0000000000000000000000000030000000000;  // -0.0000000000002274 = 0.5 * ln( 1 + -1 * 2^(-42+1) + (-1^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = -1 
assign X[4'b0011] [42] = 146'h 000000000000000000000000000C000000000;  // -0.0000000000001137 = 0.5 * ln( 1 + -1 * 2^(-43+1) + (-1^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = -1 
assign X[4'b0011] [43] = 146'h 0000000000000000000000000003000000000;  // -0.0000000000000568 = 0.5 * ln( 1 + -1 * 2^(-44+1) + (-1^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = -1 
assign X[4'b0011] [44] = 146'h 0000000000000000000000000000C00000000;  // -0.0000000000000284 = 0.5 * ln( 1 + -1 * 2^(-45+1) + (-1^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = -1 
assign X[4'b0011] [45] = 146'h 0000000000000000000000000000300000000;  // -0.0000000000000142 = 0.5 * ln( 1 + -1 * 2^(-46+1) + (-1^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = -1 
assign X[4'b0011] [46] = 146'h 00000000000000000000000000000C0000000;  // -0.0000000000000071 = 0.5 * ln( 1 + -1 * 2^(-47+1) + (-1^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = -1 
assign X[4'b0011] [47] = 146'h 0000000000000000000000000000030000000;  // -0.0000000000000036 = 0.5 * ln( 1 + -1 * 2^(-48+1) + (-1^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = -1 
assign X[4'b0011] [48] = 146'h 000000000000000000000000000000C000000;  // -0.0000000000000018 = 0.5 * ln( 1 + -1 * 2^(-49+1) + (-1^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = -1 
assign X[4'b0011] [49] = 146'h 0000000000000000000000000000003000000;  // -0.0000000000000009 = 0.5 * ln( 1 + -1 * 2^(-50+1) + (-1^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = -1 
assign X[4'b0011] [50] = 146'h 0000000000000000000000000000000C00000;  // -0.0000000000000004 = 0.5 * ln( 1 + -1 * 2^(-51+1) + (-1^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = -1 
assign X[4'b0011] [51] = 146'h 0000000000000000000000000000000300000;  // -0.0000000000000002 = 0.5 * ln( 1 + -1 * 2^(-52+1) + (-1^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = -1 
assign X[4'b0011] [52] = 146'h 00000000000000000000000000000000C0000;  // -0.0000000000000001 = 0.5 * ln( 1 + -1 * 2^(-53+1) + (-1^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = -1 
assign X[4'b0011] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-54+1) + (-1^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = -1 
assign X[4'b0011] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-55+1) + (-1^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = -1 
assign X[4'b0011] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-56+1) + (-1^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = -1 
assign X[4'b0011] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-57+1) + (-1^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = -1 
assign X[4'b0011] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-58+1) + (-1^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = -1 
assign X[4'b0011] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-59+1) + (-1^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = -1 
assign X[4'b0011] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-60+1) + (-1^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = -1 
assign X[4'b0011] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-61+1) + (-1^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = -1 
assign X[4'b0011] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-62+1) + (-1^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = -1 
assign X[4'b0011] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-63+1) + (-1^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = -1 
assign X[4'b0011] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-64+1) + (-1^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = -1 
assign X[4'b0100] [00] = 146'h 0000000430410000C03040000000000000000;  // +0.1115717756571049 = 0.5 * ln( 1 +  0 * 2^(-1+1) + ( 0^2+ 1^2) * 2^(-2*1) )   n =  1   d_n = 0+1i 
assign X[4'b0100] [01] = 146'h 0000000040300441301300000000000000000;  // +0.0303123109082174 = 0.5 * ln( 1 +  0 * 2^(-2+1) + ( 0^2+ 1^2) * 2^(-2*2) )   n =  2   d_n = 0+1i 
assign X[4'b0100] [02] = 146'h 0000000004003000444133000000000000000;  // +0.0077520932679826 = 0.5 * ln( 1 +  0 * 2^(-3+1) + ( 0^2+ 1^2) * 2^(-2*3) )   n =  3   d_n = 0+1i 
assign X[4'b0100] [03] = 146'h 0000000000400030000444400000000000000;  // +0.0019493202078287 = 0.5 * ln( 1 +  0 * 2^(-4+1) + ( 0^2+ 1^2) * 2^(-2*4) )   n =  4   d_n = 0+1i 
assign X[4'b0100] [04] = 146'h 0000000000040000300000444000000000000;  // +0.0004880429865277 = 0.5 * ln( 1 +  0 * 2^(-5+1) + ( 0^2+ 1^2) * 2^(-2*5) )   n =  5   d_n = 0+1i 
assign X[4'b0100] [05] = 146'h 0000000000004000003000000400000000000;  // +0.0001220554137636 = 0.5 * ln( 1 +  0 * 2^(-6+1) + ( 0^2+ 1^2) * 2^(-2*6) )   n =  6   d_n = 0+1i 
assign X[4'b0100] [06] = 146'h 0000000000000400000030000000000000000;  // +0.0000305166468403 = 0.5 * ln( 1 +  0 * 2^(-7+1) + ( 0^2+ 1^2) * 2^(-2*7) )   n =  7   d_n = 0+1i 
assign X[4'b0100] [07] = 146'h 0000000000000040000000300000000000000;  // +0.0000076293363242 = 0.5 * ln( 1 +  0 * 2^(-8+1) + ( 0^2+ 1^2) * 2^(-2*8) )   n =  8   d_n = 0+1i 
assign X[4'b0100] [08] = 146'h 0000000000000004000000003000000000000;  // +0.0000019073449948 = 0.5 * ln( 1 +  0 * 2^(-9+1) + ( 0^2+ 1^2) * 2^(-2*9) )   n =  9   d_n = 0+1i 
assign X[4'b0100] [09] = 146'h 0000000000000000400000000030000000000;  // +0.0000004768369308 = 0.5 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 1^2) * 2^(-2*10) )   n = 10   d_n = 0+1i 
assign X[4'b0100] [10] = 146'h 0000000000000000040000000000300000000;  // +0.0000001192092753 = 0.5 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 1^2) * 2^(-2*11) )   n = 11   d_n = 0+1i 
assign X[4'b0100] [11] = 146'h 0000000000000000004000000000003000000;  // +0.0000000298023215 = 0.5 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 1^2) * 2^(-2*12) )   n = 12   d_n = 0+1i 
assign X[4'b0100] [12] = 146'h 0000000000000000000400000000000000000;  // +0.0000000074505806 = 0.5 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 1^2) * 2^(-2*13) )   n = 13   d_n = 0+1i 
assign X[4'b0100] [13] = 146'h 0000000000000000000040000000000000000;  // +0.0000000018626451 = 0.5 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 1^2) * 2^(-2*14) )   n = 14   d_n = 0+1i 
assign X[4'b0100] [14] = 146'h 0000000000000000000004000000000000000;  // +0.0000000004656613 = 0.5 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 1^2) * 2^(-2*15) )   n = 15   d_n = 0+1i 
assign X[4'b0100] [15] = 146'h 0000000000000000000000400000000000000;  // +0.0000000001164153 = 0.5 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 1^2) * 2^(-2*16) )   n = 16   d_n = 0+1i 
assign X[4'b0100] [16] = 146'h 0000000000000000000000040000000000000;  // +0.0000000000291038 = 0.5 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 1^2) * 2^(-2*17) )   n = 17   d_n = 0+1i 
assign X[4'b0100] [17] = 146'h 0000000000000000000000004000000000000;  // +0.0000000000072760 = 0.5 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 1^2) * 2^(-2*18) )   n = 18   d_n = 0+1i 
assign X[4'b0100] [18] = 146'h 0000000000000000000000000400000000000;  // +0.0000000000018190 = 0.5 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 1^2) * 2^(-2*19) )   n = 19   d_n = 0+1i 
assign X[4'b0100] [19] = 146'h 0000000000000000000000000040000000000;  // +0.0000000000004547 = 0.5 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 1^2) * 2^(-2*20) )   n = 20   d_n = 0+1i 
assign X[4'b0100] [20] = 146'h 0000000000000000000000000004000000000;  // +0.0000000000001137 = 0.5 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 1^2) * 2^(-2*21) )   n = 21   d_n = 0+1i 
assign X[4'b0100] [21] = 146'h 0000000000000000000000000000400000000;  // +0.0000000000000284 = 0.5 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 1^2) * 2^(-2*22) )   n = 22   d_n = 0+1i 
assign X[4'b0100] [22] = 146'h 0000000000000000000000000000040000000;  // +0.0000000000000071 = 0.5 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 1^2) * 2^(-2*23) )   n = 23   d_n = 0+1i 
assign X[4'b0100] [23] = 146'h 0000000000000000000000000000004000000;  // +0.0000000000000018 = 0.5 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 1^2) * 2^(-2*24) )   n = 24   d_n = 0+1i 
assign X[4'b0100] [24] = 146'h 0000000000000000000000000000000400000;  // +0.0000000000000004 = 0.5 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 1^2) * 2^(-2*25) )   n = 25   d_n = 0+1i 
assign X[4'b0100] [25] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 1^2) * 2^(-2*26) )   n = 26   d_n = 0+1i 
assign X[4'b0100] [26] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 1^2) * 2^(-2*27) )   n = 27   d_n = 0+1i 
assign X[4'b0100] [27] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 1^2) * 2^(-2*28) )   n = 28   d_n = 0+1i 
assign X[4'b0100] [28] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 1^2) * 2^(-2*29) )   n = 29   d_n = 0+1i 
assign X[4'b0100] [29] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 1^2) * 2^(-2*30) )   n = 30   d_n = 0+1i 
assign X[4'b0100] [30] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 1^2) * 2^(-2*31) )   n = 31   d_n = 0+1i 
assign X[4'b0100] [31] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 1^2) * 2^(-2*32) )   n = 32   d_n = 0+1i 
assign X[4'b0100] [32] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 1^2) * 2^(-2*33) )   n = 33   d_n = 0+1i 
assign X[4'b0100] [33] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 1^2) * 2^(-2*34) )   n = 34   d_n = 0+1i 
assign X[4'b0100] [34] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 1^2) * 2^(-2*35) )   n = 35   d_n = 0+1i 
assign X[4'b0100] [35] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 1^2) * 2^(-2*36) )   n = 36   d_n = 0+1i 
assign X[4'b0100] [36] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 1^2) * 2^(-2*37) )   n = 37   d_n = 0+1i 
assign X[4'b0100] [37] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 1^2) * 2^(-2*38) )   n = 38   d_n = 0+1i 
assign X[4'b0100] [38] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 1^2) * 2^(-2*39) )   n = 39   d_n = 0+1i 
assign X[4'b0100] [39] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 1^2) * 2^(-2*40) )   n = 40   d_n = 0+1i 
assign X[4'b0100] [40] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 1^2) * 2^(-2*41) )   n = 41   d_n = 0+1i 
assign X[4'b0100] [41] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 1^2) * 2^(-2*42) )   n = 42   d_n = 0+1i 
assign X[4'b0100] [42] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 1^2) * 2^(-2*43) )   n = 43   d_n = 0+1i 
assign X[4'b0100] [43] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 1^2) * 2^(-2*44) )   n = 44   d_n = 0+1i 
assign X[4'b0100] [44] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 1^2) * 2^(-2*45) )   n = 45   d_n = 0+1i 
assign X[4'b0100] [45] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 1^2) * 2^(-2*46) )   n = 46   d_n = 0+1i 
assign X[4'b0100] [46] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 1^2) * 2^(-2*47) )   n = 47   d_n = 0+1i 
assign X[4'b0100] [47] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 1^2) * 2^(-2*48) )   n = 48   d_n = 0+1i 
assign X[4'b0100] [48] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 1^2) * 2^(-2*49) )   n = 49   d_n = 0+1i 
assign X[4'b0100] [49] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 1^2) * 2^(-2*50) )   n = 50   d_n = 0+1i 
assign X[4'b0100] [50] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 1^2) * 2^(-2*51) )   n = 51   d_n = 0+1i 
assign X[4'b0100] [51] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 1^2) * 2^(-2*52) )   n = 52   d_n = 0+1i 
assign X[4'b0100] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 1^2) * 2^(-2*53) )   n = 53   d_n = 0+1i 
assign X[4'b0100] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 1^2) * 2^(-2*54) )   n = 54   d_n = 0+1i 
assign X[4'b0100] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 1^2) * 2^(-2*55) )   n = 55   d_n = 0+1i 
assign X[4'b0100] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 1^2) * 2^(-2*56) )   n = 56   d_n = 0+1i 
assign X[4'b0100] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 1^2) * 2^(-2*57) )   n = 57   d_n = 0+1i 
assign X[4'b0100] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 1^2) * 2^(-2*58) )   n = 58   d_n = 0+1i 
assign X[4'b0100] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 1^2) * 2^(-2*59) )   n = 59   d_n = 0+1i 
assign X[4'b0100] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 1^2) * 2^(-2*60) )   n = 60   d_n = 0+1i 
assign X[4'b0100] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 1^2) * 2^(-2*61) )   n = 61   d_n = 0+1i 
assign X[4'b0100] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 1^2) * 2^(-2*62) )   n = 62   d_n = 0+1i 
assign X[4'b0100] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 1^2) * 2^(-2*63) )   n = 63   d_n = 0+1i 
assign X[4'b0100] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 1^2) * 2^(-2*64) )   n = 64   d_n = 0+1i 
assign X[4'b0101] [00] = 146'h 0000004311104100103000000000000000000;  // +0.4581453659370776 = 0.5 * ln( 1 +  1 * 2^(-1+1) + ( 1^2+ 1^2) * 2^(-2*1) )   n =  1   d_n = 1+1i 
assign X[4'b0101] [01] = 146'h 000000100C041104033000000000000000000;  // +0.2427539078908503 = 0.5 * ln( 1 +  1 * 2^(-2+1) + ( 1^2+ 1^2) * 2^(-2*2) )   n =  2   d_n = 1+1i 
assign X[4'b0101] [02] = 146'h 000000040030C104C04300000000000000000;  // +0.1239180819522907 = 0.5 * ln( 1 +  1 * 2^(-3+1) + ( 1^2+ 1^2) * 2^(-2*3) )   n =  3   d_n = 1+1i 
assign X[4'b0101] [03] = 146'h 000000010000CC104044C0000000000000000;  // +0.0623517392504787 = 0.5 * ln( 1 +  1 * 2^(-4+1) + ( 1^2+ 1^2) * 2^(-2*4) )   n =  4   d_n = 1+1i 
assign X[4'b0101] [04] = 146'h 0000000040000330C41010000000000000000;  // +0.0312305848118681 = 0.5 * ln( 1 +  1 * 2^(-5+1) + ( 1^2+ 1^2) * 2^(-2*5) )   n =  5   d_n = 1+1i 
assign X[4'b0101] [05] = 146'h 000000001000000CCC1104000000000000000;  // +0.0156225157283291 = 0.5 * ln( 1 +  1 * 2^(-6+1) + ( 1^2+ 1^2) * 2^(-2*6) )   n =  6   d_n = 1+1i 
assign X[4'b0101] [06] = 146'h 00000000040000003330C4400000000000000;  // +0.0078121858105703 = 0.5 * ln( 1 +  1 * 2^(-7+1) + ( 1^2+ 1^2) * 2^(-2*7) )   n =  7   d_n = 1+1i 
assign X[4'b0101] [07] = 146'h 000000000100000000CCCC100000000000000;  // +0.0039062104956732 = 0.5 * ln( 1 +  1 * 2^(-8+1) + ( 1^2+ 1^2) * 2^(-2*8) )   n =  8   d_n = 1+1i 
assign X[4'b0101] [08] = 146'h 0000000000400000000333300000000000000;  // +0.0019531200474755 = 0.5 * ln( 1 +  1 * 2^(-9+1) + ( 1^2+ 1^2) * 2^(-2*9) )   n =  9   d_n = 1+1i 
assign X[4'b0101] [09] = 146'h 000000000010000000000CCD0000000000000;  // +0.0009765618800270 = 0.5 * ln( 1 +  1 * 2^(-10+1) + ( 1^2+ 1^2) * 2^(-2*10) )   n = 10   d_n = 1+1i 
assign X[4'b0101] [10] = 146'h 0000000000040000000000334000000000000;  // +0.0004882811724466 = 0.5 * ln( 1 +  1 * 2^(-11+1) + ( 1^2+ 1^2) * 2^(-2*11) )   n = 11   d_n = 1+1i 
assign X[4'b0101] [11] = 146'h 000000000001000000000000D000000000000;  // +0.0002441406153023 = 0.5 * ln( 1 +  1 * 2^(-12+1) + ( 1^2+ 1^2) * 2^(-2*12) )   n = 12   d_n = 1+1i 
assign X[4'b0101] [12] = 146'h 0000000000004000000000000400000000000;  // +0.0001220703112875 = 0.5 * ln( 1 +  1 * 2^(-13+1) + ( 1^2+ 1^2) * 2^(-2*13) )   n = 13   d_n = 1+1i 
assign X[4'b0101] [13] = 146'h 0000000000001000000000000000000000000;  // +0.0000610351560984 = 0.5 * ln( 1 +  1 * 2^(-14+1) + ( 1^2+ 1^2) * 2^(-2*14) )   n = 14   d_n = 1+1i 
assign X[4'b0101] [14] = 146'h 0000000000000400000000000000000000000;  // +0.0000305175781061 = 0.5 * ln( 1 +  1 * 2^(-15+1) + ( 1^2+ 1^2) * 2^(-2*15) )   n = 15   d_n = 1+1i 
assign X[4'b0101] [15] = 146'h 0000000000000100000000000000000000000;  // +0.0000152587890601 = 0.5 * ln( 1 +  1 * 2^(-16+1) + ( 1^2+ 1^2) * 2^(-2*16) )   n = 16   d_n = 1+1i 
assign X[4'b0101] [16] = 146'h 0000000000000040000000000000000000000;  // +0.0000076293945310 = 0.5 * ln( 1 +  1 * 2^(-17+1) + ( 1^2+ 1^2) * 2^(-2*17) )   n = 17   d_n = 1+1i 
assign X[4'b0101] [17] = 146'h 0000000000000010000000000000000000000;  // +0.0000038146972656 = 0.5 * ln( 1 +  1 * 2^(-18+1) + ( 1^2+ 1^2) * 2^(-2*18) )   n = 18   d_n = 1+1i 
assign X[4'b0101] [18] = 146'h 0000000000000004000000000000000000000;  // +0.0000019073486328 = 0.5 * ln( 1 +  1 * 2^(-19+1) + ( 1^2+ 1^2) * 2^(-2*19) )   n = 19   d_n = 1+1i 
assign X[4'b0101] [19] = 146'h 0000000000000001000000000000000000000;  // +0.0000009536743164 = 0.5 * ln( 1 +  1 * 2^(-20+1) + ( 1^2+ 1^2) * 2^(-2*20) )   n = 20   d_n = 1+1i 
assign X[4'b0101] [20] = 146'h 0000000000000000400000000000000000000;  // +0.0000004768371582 = 0.5 * ln( 1 +  1 * 2^(-21+1) + ( 1^2+ 1^2) * 2^(-2*21) )   n = 21   d_n = 1+1i 
assign X[4'b0101] [21] = 146'h 0000000000000000100000000000000000000;  // +0.0000002384185791 = 0.5 * ln( 1 +  1 * 2^(-22+1) + ( 1^2+ 1^2) * 2^(-2*22) )   n = 22   d_n = 1+1i 
assign X[4'b0101] [22] = 146'h 0000000000000000040000000000000000000;  // +0.0000001192092896 = 0.5 * ln( 1 +  1 * 2^(-23+1) + ( 1^2+ 1^2) * 2^(-2*23) )   n = 23   d_n = 1+1i 
assign X[4'b0101] [23] = 146'h 0000000000000000010000000000000000000;  // +0.0000000596046448 = 0.5 * ln( 1 +  1 * 2^(-24+1) + ( 1^2+ 1^2) * 2^(-2*24) )   n = 24   d_n = 1+1i 
assign X[4'b0101] [24] = 146'h 0000000000000000004000000000000000000;  // +0.0000000298023224 = 0.5 * ln( 1 +  1 * 2^(-25+1) + ( 1^2+ 1^2) * 2^(-2*25) )   n = 25   d_n = 1+1i 
assign X[4'b0101] [25] = 146'h 0000000000000000001000000000000100000;  // +0.0000000149011611 = 0.5 * ln( 1 +  1 * 2^(-26+1) + ( 1^2+ 1^2) * 2^(-2*26) )   n = 26   d_n = 1+1i 
assign X[4'b0101] [26] = 146'h 0000000000000000000400000000000000000;  // +0.0000000074505806 = 0.5 * ln( 1 +  1 * 2^(-27+1) + ( 1^2+ 1^2) * 2^(-2*27) )   n = 27   d_n = 1+1i 
assign X[4'b0101] [27] = 146'h 0000000000000000000100000000000000000;  // +0.0000000037252903 = 0.5 * ln( 1 +  1 * 2^(-28+1) + ( 1^2+ 1^2) * 2^(-2*28) )   n = 28   d_n = 1+1i 
assign X[4'b0101] [28] = 146'h 0000000000000000000040000000000000000;  // +0.0000000018626451 = 0.5 * ln( 1 +  1 * 2^(-29+1) + ( 1^2+ 1^2) * 2^(-2*29) )   n = 29   d_n = 1+1i 
assign X[4'b0101] [29] = 146'h 0000000000000000000010000000000000000;  // +0.0000000009313226 = 0.5 * ln( 1 +  1 * 2^(-30+1) + ( 1^2+ 1^2) * 2^(-2*30) )   n = 30   d_n = 1+1i 
assign X[4'b0101] [30] = 146'h 0000000000000000000004000000000000000;  // +0.0000000004656613 = 0.5 * ln( 1 +  1 * 2^(-31+1) + ( 1^2+ 1^2) * 2^(-2*31) )   n = 31   d_n = 1+1i 
assign X[4'b0101] [31] = 146'h 0000000000000000000001000000000000000;  // +0.0000000002328306 = 0.5 * ln( 1 +  1 * 2^(-32+1) + ( 1^2+ 1^2) * 2^(-2*32) )   n = 32   d_n = 1+1i 
assign X[4'b0101] [32] = 146'h 0000000000000000000000400000000000000;  // +0.0000000001164153 = 0.5 * ln( 1 +  1 * 2^(-33+1) + ( 1^2+ 1^2) * 2^(-2*33) )   n = 33   d_n = 1+1i 
assign X[4'b0101] [33] = 146'h 0000000000000000000000100000000000000;  // +0.0000000000582077 = 0.5 * ln( 1 +  1 * 2^(-34+1) + ( 1^2+ 1^2) * 2^(-2*34) )   n = 34   d_n = 1+1i 
assign X[4'b0101] [34] = 146'h 0000000000000000000000040000000000000;  // +0.0000000000291038 = 0.5 * ln( 1 +  1 * 2^(-35+1) + ( 1^2+ 1^2) * 2^(-2*35) )   n = 35   d_n = 1+1i 
assign X[4'b0101] [35] = 146'h 0000000000000000000000010000000000000;  // +0.0000000000145519 = 0.5 * ln( 1 +  1 * 2^(-36+1) + ( 1^2+ 1^2) * 2^(-2*36) )   n = 36   d_n = 1+1i 
assign X[4'b0101] [36] = 146'h 0000000000000000000000004000000000000;  // +0.0000000000072760 = 0.5 * ln( 1 +  1 * 2^(-37+1) + ( 1^2+ 1^2) * 2^(-2*37) )   n = 37   d_n = 1+1i 
assign X[4'b0101] [37] = 146'h 0000000000000000000000001000000000000;  // +0.0000000000036380 = 0.5 * ln( 1 +  1 * 2^(-38+1) + ( 1^2+ 1^2) * 2^(-2*38) )   n = 38   d_n = 1+1i 
assign X[4'b0101] [38] = 146'h 0000000000000000000000000400000000000;  // +0.0000000000018190 = 0.5 * ln( 1 +  1 * 2^(-39+1) + ( 1^2+ 1^2) * 2^(-2*39) )   n = 39   d_n = 1+1i 
assign X[4'b0101] [39] = 146'h 0000000000000000000000000100000000000;  // +0.0000000000009095 = 0.5 * ln( 1 +  1 * 2^(-40+1) + ( 1^2+ 1^2) * 2^(-2*40) )   n = 40   d_n = 1+1i 
assign X[4'b0101] [40] = 146'h 0000000000000000000000000040000000000;  // +0.0000000000004547 = 0.5 * ln( 1 +  1 * 2^(-41+1) + ( 1^2+ 1^2) * 2^(-2*41) )   n = 41   d_n = 1+1i 
assign X[4'b0101] [41] = 146'h 0000000000000000000000000010000000000;  // +0.0000000000002274 = 0.5 * ln( 1 +  1 * 2^(-42+1) + ( 1^2+ 1^2) * 2^(-2*42) )   n = 42   d_n = 1+1i 
assign X[4'b0101] [42] = 146'h 0000000000000000000000000004000000000;  // +0.0000000000001137 = 0.5 * ln( 1 +  1 * 2^(-43+1) + ( 1^2+ 1^2) * 2^(-2*43) )   n = 43   d_n = 1+1i 
assign X[4'b0101] [43] = 146'h 0000000000000000000000000001000000000;  // +0.0000000000000568 = 0.5 * ln( 1 +  1 * 2^(-44+1) + ( 1^2+ 1^2) * 2^(-2*44) )   n = 44   d_n = 1+1i 
assign X[4'b0101] [44] = 146'h 0000000000000000000000000000400000000;  // +0.0000000000000284 = 0.5 * ln( 1 +  1 * 2^(-45+1) + ( 1^2+ 1^2) * 2^(-2*45) )   n = 45   d_n = 1+1i 
assign X[4'b0101] [45] = 146'h 0000000000000000000000000000100000000;  // +0.0000000000000142 = 0.5 * ln( 1 +  1 * 2^(-46+1) + ( 1^2+ 1^2) * 2^(-2*46) )   n = 46   d_n = 1+1i 
assign X[4'b0101] [46] = 146'h 0000000000000000000000000000040000000;  // +0.0000000000000071 = 0.5 * ln( 1 +  1 * 2^(-47+1) + ( 1^2+ 1^2) * 2^(-2*47) )   n = 47   d_n = 1+1i 
assign X[4'b0101] [47] = 146'h 0000000000000000000000000000010000000;  // +0.0000000000000036 = 0.5 * ln( 1 +  1 * 2^(-48+1) + ( 1^2+ 1^2) * 2^(-2*48) )   n = 48   d_n = 1+1i 
assign X[4'b0101] [48] = 146'h 0000000000000000000000000000004000000;  // +0.0000000000000018 = 0.5 * ln( 1 +  1 * 2^(-49+1) + ( 1^2+ 1^2) * 2^(-2*49) )   n = 49   d_n = 1+1i 
assign X[4'b0101] [49] = 146'h 0000000000000000000000000000001000000;  // +0.0000000000000009 = 0.5 * ln( 1 +  1 * 2^(-50+1) + ( 1^2+ 1^2) * 2^(-2*50) )   n = 50   d_n = 1+1i 
assign X[4'b0101] [50] = 146'h 0000000000000000000000000000000400000;  // +0.0000000000000004 = 0.5 * ln( 1 +  1 * 2^(-51+1) + ( 1^2+ 1^2) * 2^(-2*51) )   n = 51   d_n = 1+1i 
assign X[4'b0101] [51] = 146'h 0000000000000000000000000000000100000;  // +0.0000000000000002 = 0.5 * ln( 1 +  1 * 2^(-52+1) + ( 1^2+ 1^2) * 2^(-2*52) )   n = 52   d_n = 1+1i 
assign X[4'b0101] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-53+1) + ( 1^2+ 1^2) * 2^(-2*53) )   n = 53   d_n = 1+1i 
assign X[4'b0101] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-54+1) + ( 1^2+ 1^2) * 2^(-2*54) )   n = 54   d_n = 1+1i 
assign X[4'b0101] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-55+1) + ( 1^2+ 1^2) * 2^(-2*55) )   n = 55   d_n = 1+1i 
assign X[4'b0101] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-56+1) + ( 1^2+ 1^2) * 2^(-2*56) )   n = 56   d_n = 1+1i 
assign X[4'b0101] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-57+1) + ( 1^2+ 1^2) * 2^(-2*57) )   n = 57   d_n = 1+1i 
assign X[4'b0101] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-58+1) + ( 1^2+ 1^2) * 2^(-2*58) )   n = 58   d_n = 1+1i 
assign X[4'b0101] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-59+1) + ( 1^2+ 1^2) * 2^(-2*59) )   n = 59   d_n = 1+1i 
assign X[4'b0101] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-60+1) + ( 1^2+ 1^2) * 2^(-2*60) )   n = 60   d_n = 1+1i 
assign X[4'b0101] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-61+1) + ( 1^2+ 1^2) * 2^(-2*61) )   n = 61   d_n = 1+1i 
assign X[4'b0101] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-62+1) + ( 1^2+ 1^2) * 2^(-2*62) )   n = 62   d_n = 1+1i 
assign X[4'b0101] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-63+1) + ( 1^2+ 1^2) * 2^(-2*63) )   n = 63   d_n = 1+1i 
assign X[4'b0101] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-64+1) + ( 1^2+ 1^2) * 2^(-2*64) )   n = 64   d_n = 1+1i 
assign X[4'b0110] [00] = 146'h 0000000430410000C03040000000000000000;  // +0.1115717756571049 = 0.5 * ln( 1 +  0 * 2^(-1+1) + ( 0^2+ 1^2) * 2^(-2*1) )   n =  1   d_n = 0+1i 
assign X[4'b0110] [01] = 146'h 0000000040300441301300000000000000000;  // +0.0303123109082174 = 0.5 * ln( 1 +  0 * 2^(-2+1) + ( 0^2+ 1^2) * 2^(-2*2) )   n =  2   d_n = 0+1i 
assign X[4'b0110] [02] = 146'h 0000000004003000444133000000000000000;  // +0.0077520932679826 = 0.5 * ln( 1 +  0 * 2^(-3+1) + ( 0^2+ 1^2) * 2^(-2*3) )   n =  3   d_n = 0+1i 
assign X[4'b0110] [03] = 146'h 0000000000400030000444400000000000000;  // +0.0019493202078287 = 0.5 * ln( 1 +  0 * 2^(-4+1) + ( 0^2+ 1^2) * 2^(-2*4) )   n =  4   d_n = 0+1i 
assign X[4'b0110] [04] = 146'h 0000000000040000300000444000000000000;  // +0.0004880429865277 = 0.5 * ln( 1 +  0 * 2^(-5+1) + ( 0^2+ 1^2) * 2^(-2*5) )   n =  5   d_n = 0+1i 
assign X[4'b0110] [05] = 146'h 0000000000004000003000000400000000000;  // +0.0001220554137636 = 0.5 * ln( 1 +  0 * 2^(-6+1) + ( 0^2+ 1^2) * 2^(-2*6) )   n =  6   d_n = 0+1i 
assign X[4'b0110] [06] = 146'h 0000000000000400000030000000000000000;  // +0.0000305166468403 = 0.5 * ln( 1 +  0 * 2^(-7+1) + ( 0^2+ 1^2) * 2^(-2*7) )   n =  7   d_n = 0+1i 
assign X[4'b0110] [07] = 146'h 0000000000000040000000300000000000000;  // +0.0000076293363242 = 0.5 * ln( 1 +  0 * 2^(-8+1) + ( 0^2+ 1^2) * 2^(-2*8) )   n =  8   d_n = 0+1i 
assign X[4'b0110] [08] = 146'h 0000000000000004000000003000000000000;  // +0.0000019073449948 = 0.5 * ln( 1 +  0 * 2^(-9+1) + ( 0^2+ 1^2) * 2^(-2*9) )   n =  9   d_n = 0+1i 
assign X[4'b0110] [09] = 146'h 0000000000000000400000000030000000000;  // +0.0000004768369308 = 0.5 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 1^2) * 2^(-2*10) )   n = 10   d_n = 0+1i 
assign X[4'b0110] [10] = 146'h 0000000000000000040000000000300000000;  // +0.0000001192092753 = 0.5 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 1^2) * 2^(-2*11) )   n = 11   d_n = 0+1i 
assign X[4'b0110] [11] = 146'h 0000000000000000004000000000003000000;  // +0.0000000298023215 = 0.5 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 1^2) * 2^(-2*12) )   n = 12   d_n = 0+1i 
assign X[4'b0110] [12] = 146'h 0000000000000000000400000000000000000;  // +0.0000000074505806 = 0.5 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 1^2) * 2^(-2*13) )   n = 13   d_n = 0+1i 
assign X[4'b0110] [13] = 146'h 0000000000000000000040000000000000000;  // +0.0000000018626451 = 0.5 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 1^2) * 2^(-2*14) )   n = 14   d_n = 0+1i 
assign X[4'b0110] [14] = 146'h 0000000000000000000004000000000000000;  // +0.0000000004656613 = 0.5 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 1^2) * 2^(-2*15) )   n = 15   d_n = 0+1i 
assign X[4'b0110] [15] = 146'h 0000000000000000000000400000000000000;  // +0.0000000001164153 = 0.5 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 1^2) * 2^(-2*16) )   n = 16   d_n = 0+1i 
assign X[4'b0110] [16] = 146'h 0000000000000000000000040000000000000;  // +0.0000000000291038 = 0.5 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 1^2) * 2^(-2*17) )   n = 17   d_n = 0+1i 
assign X[4'b0110] [17] = 146'h 0000000000000000000000004000000000000;  // +0.0000000000072760 = 0.5 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 1^2) * 2^(-2*18) )   n = 18   d_n = 0+1i 
assign X[4'b0110] [18] = 146'h 0000000000000000000000000400000000000;  // +0.0000000000018190 = 0.5 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 1^2) * 2^(-2*19) )   n = 19   d_n = 0+1i 
assign X[4'b0110] [19] = 146'h 0000000000000000000000000040000000000;  // +0.0000000000004547 = 0.5 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 1^2) * 2^(-2*20) )   n = 20   d_n = 0+1i 
assign X[4'b0110] [20] = 146'h 0000000000000000000000000004000000000;  // +0.0000000000001137 = 0.5 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 1^2) * 2^(-2*21) )   n = 21   d_n = 0+1i 
assign X[4'b0110] [21] = 146'h 0000000000000000000000000000400000000;  // +0.0000000000000284 = 0.5 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 1^2) * 2^(-2*22) )   n = 22   d_n = 0+1i 
assign X[4'b0110] [22] = 146'h 0000000000000000000000000000040000000;  // +0.0000000000000071 = 0.5 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 1^2) * 2^(-2*23) )   n = 23   d_n = 0+1i 
assign X[4'b0110] [23] = 146'h 0000000000000000000000000000004000000;  // +0.0000000000000018 = 0.5 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 1^2) * 2^(-2*24) )   n = 24   d_n = 0+1i 
assign X[4'b0110] [24] = 146'h 0000000000000000000000000000000400000;  // +0.0000000000000004 = 0.5 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 1^2) * 2^(-2*25) )   n = 25   d_n = 0+1i 
assign X[4'b0110] [25] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 1^2) * 2^(-2*26) )   n = 26   d_n = 0+1i 
assign X[4'b0110] [26] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 1^2) * 2^(-2*27) )   n = 27   d_n = 0+1i 
assign X[4'b0110] [27] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 1^2) * 2^(-2*28) )   n = 28   d_n = 0+1i 
assign X[4'b0110] [28] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 1^2) * 2^(-2*29) )   n = 29   d_n = 0+1i 
assign X[4'b0110] [29] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 1^2) * 2^(-2*30) )   n = 30   d_n = 0+1i 
assign X[4'b0110] [30] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 1^2) * 2^(-2*31) )   n = 31   d_n = 0+1i 
assign X[4'b0110] [31] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 1^2) * 2^(-2*32) )   n = 32   d_n = 0+1i 
assign X[4'b0110] [32] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 1^2) * 2^(-2*33) )   n = 33   d_n = 0+1i 
assign X[4'b0110] [33] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 1^2) * 2^(-2*34) )   n = 34   d_n = 0+1i 
assign X[4'b0110] [34] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 1^2) * 2^(-2*35) )   n = 35   d_n = 0+1i 
assign X[4'b0110] [35] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 1^2) * 2^(-2*36) )   n = 36   d_n = 0+1i 
assign X[4'b0110] [36] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 1^2) * 2^(-2*37) )   n = 37   d_n = 0+1i 
assign X[4'b0110] [37] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 1^2) * 2^(-2*38) )   n = 38   d_n = 0+1i 
assign X[4'b0110] [38] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 1^2) * 2^(-2*39) )   n = 39   d_n = 0+1i 
assign X[4'b0110] [39] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 1^2) * 2^(-2*40) )   n = 40   d_n = 0+1i 
assign X[4'b0110] [40] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 1^2) * 2^(-2*41) )   n = 41   d_n = 0+1i 
assign X[4'b0110] [41] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 1^2) * 2^(-2*42) )   n = 42   d_n = 0+1i 
assign X[4'b0110] [42] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 1^2) * 2^(-2*43) )   n = 43   d_n = 0+1i 
assign X[4'b0110] [43] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 1^2) * 2^(-2*44) )   n = 44   d_n = 0+1i 
assign X[4'b0110] [44] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 1^2) * 2^(-2*45) )   n = 45   d_n = 0+1i 
assign X[4'b0110] [45] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 1^2) * 2^(-2*46) )   n = 46   d_n = 0+1i 
assign X[4'b0110] [46] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 1^2) * 2^(-2*47) )   n = 47   d_n = 0+1i 
assign X[4'b0110] [47] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 1^2) * 2^(-2*48) )   n = 48   d_n = 0+1i 
assign X[4'b0110] [48] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 1^2) * 2^(-2*49) )   n = 49   d_n = 0+1i 
assign X[4'b0110] [49] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 1^2) * 2^(-2*50) )   n = 50   d_n = 0+1i 
assign X[4'b0110] [50] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 1^2) * 2^(-2*51) )   n = 51   d_n = 0+1i 
assign X[4'b0110] [51] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 1^2) * 2^(-2*52) )   n = 52   d_n = 0+1i 
assign X[4'b0110] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 1^2) * 2^(-2*53) )   n = 53   d_n = 0+1i 
assign X[4'b0110] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 1^2) * 2^(-2*54) )   n = 54   d_n = 0+1i 
assign X[4'b0110] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 1^2) * 2^(-2*55) )   n = 55   d_n = 0+1i 
assign X[4'b0110] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 1^2) * 2^(-2*56) )   n = 56   d_n = 0+1i 
assign X[4'b0110] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 1^2) * 2^(-2*57) )   n = 57   d_n = 0+1i 
assign X[4'b0110] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 1^2) * 2^(-2*58) )   n = 58   d_n = 0+1i 
assign X[4'b0110] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 1^2) * 2^(-2*59) )   n = 59   d_n = 0+1i 
assign X[4'b0110] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 1^2) * 2^(-2*60) )   n = 60   d_n = 0+1i 
assign X[4'b0110] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 1^2) * 2^(-2*61) )   n = 61   d_n = 0+1i 
assign X[4'b0110] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 1^2) * 2^(-2*62) )   n = 62   d_n = 0+1i 
assign X[4'b0110] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 1^2) * 2^(-2*63) )   n = 63   d_n = 0+1i 
assign X[4'b0110] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 1^2) * 2^(-2*64) )   n = 64   d_n = 0+1i 
assign X[4'b0111] [00] = 146'h 000000C443104303100000000000000000000;  // -0.3465735902799726 = 0.5 * ln( 1 + -1 * 2^(-1+1) + (-1^2+ 1^2) * 2^(-2*1) )   n =  1   d_n = -1+1i 
assign X[4'b0111] [01] = 146'h 00000030100CC303303200000000000000000;  // -0.2350018146228677 = 0.5 * ln( 1 + -1 * 2^(-2+1) + (-1^2+ 1^2) * 2^(-2*2) )   n =  2   d_n = -1+1i 
assign X[4'b0111] [02] = 146'h 0000000C004C430C10C100000000000000000;  // -0.1234300389657629 = 0.5 * ln( 1 + -1 * 2^(-3+1) + (-1^2+ 1^2) * 2^(-2*3) )   n =  3   d_n = -1+1i 
assign X[4'b0111] [03] = 146'h 0000000300013030C0CC20000000000000000;  // -0.0623212226036383 = 0.5 * ln( 1 + -1 * 2^(-4+1) + (-1^2+ 1^2) * 2^(-2*4) )   n =  4   d_n = -1+1i 
assign X[4'b0111] [04] = 146'h 00000000C00004CC4C3030000000000000000;  // -0.0312286774668733 = 0.5 * ln( 1 + -1 * 2^(-5+1) + (-1^2+ 1^2) * 2^(-2*5) )   n =  5   d_n = -1+1i 
assign X[4'b0111] [05] = 146'h 000000003000001330330C000000000000000;  // -0.0156223965190538 = 0.5 * ln( 1 + -1 * 2^(-6+1) + (-1^2+ 1^2) * 2^(-2*6) )   n =  6   d_n = -1+1i 
assign X[4'b0111] [06] = 146'h 000000000C0000004CCC4D000000000000000;  // -0.0078121783599899 = 0.5 * ln( 1 + -1 * 2^(-7+1) + (-1^2+ 1^2) * 2^(-2*7) )   n =  7   d_n = -1+1i 
assign X[4'b0111] [07] = 146'h 0000000003000000013330400000000000000;  // -0.0039062100300119 = 0.5 * ln( 1 + -1 * 2^(-8+1) + (-1^2+ 1^2) * 2^(-2*8) )   n =  8   d_n = -1+1i 
assign X[4'b0111] [08] = 146'h 0000000000C000000004CCD00000000000000;  // -0.0019531200183716 = 0.5 * ln( 1 + -1 * 2^(-9+1) + (-1^2+ 1^2) * 2^(-2*9) )   n =  9   d_n = -1+1i 
assign X[4'b0111] [09] = 146'h 0000000000300000000013340000000000000;  // -0.0009765618782081 = 0.5 * ln( 1 + -1 * 2^(-10+1) + (-1^2+ 1^2) * 2^(-2*10) )   n = 10   d_n = -1+1i 
assign X[4'b0111] [10] = 146'h 00000000000C00000000004D0000000000000;  // -0.0004882811723329 = 0.5 * ln( 1 + -1 * 2^(-11+1) + (-1^2+ 1^2) * 2^(-2*11) )   n = 11   d_n = -1+1i 
assign X[4'b0111] [11] = 146'h 0000000000030000000000014000000000000;  // -0.0002441406152952 = 0.5 * ln( 1 + -1 * 2^(-12+1) + (-1^2+ 1^2) * 2^(-2*12) )   n = 12   d_n = -1+1i 
assign X[4'b0111] [12] = 146'h 000000000000C000000000000800000000000;  // -0.0001220703112871 = 0.5 * ln( 1 + -1 * 2^(-13+1) + (-1^2+ 1^2) * 2^(-2*13) )   n = 13   d_n = -1+1i 
assign X[4'b0111] [13] = 146'h 0000000000003000000000000000000000000;  // -0.0000610351560984 = 0.5 * ln( 1 + -1 * 2^(-14+1) + (-1^2+ 1^2) * 2^(-2*14) )   n = 14   d_n = -1+1i 
assign X[4'b0111] [14] = 146'h 0000000000000C00000000000000000000000;  // -0.0000305175781061 = 0.5 * ln( 1 + -1 * 2^(-15+1) + (-1^2+ 1^2) * 2^(-2*15) )   n = 15   d_n = -1+1i 
assign X[4'b0111] [15] = 146'h 0000000000000300000000000000000000000;  // -0.0000152587890601 = 0.5 * ln( 1 + -1 * 2^(-16+1) + (-1^2+ 1^2) * 2^(-2*16) )   n = 16   d_n = -1+1i 
assign X[4'b0111] [16] = 146'h 00000000000000C0000000000000000000000;  // -0.0000076293945310 = 0.5 * ln( 1 + -1 * 2^(-17+1) + (-1^2+ 1^2) * 2^(-2*17) )   n = 17   d_n = -1+1i 
assign X[4'b0111] [17] = 146'h 0000000000000030000000000000000000000;  // -0.0000038146972656 = 0.5 * ln( 1 + -1 * 2^(-18+1) + (-1^2+ 1^2) * 2^(-2*18) )   n = 18   d_n = -1+1i 
assign X[4'b0111] [18] = 146'h 000000000000000C000000000000000000000;  // -0.0000019073486328 = 0.5 * ln( 1 + -1 * 2^(-19+1) + (-1^2+ 1^2) * 2^(-2*19) )   n = 19   d_n = -1+1i 
assign X[4'b0111] [19] = 146'h 0000000000000003000000000000000000000;  // -0.0000009536743164 = 0.5 * ln( 1 + -1 * 2^(-20+1) + (-1^2+ 1^2) * 2^(-2*20) )   n = 20   d_n = -1+1i 
assign X[4'b0111] [20] = 146'h 0000000000000000C00000000000000000000;  // -0.0000004768371582 = 0.5 * ln( 1 + -1 * 2^(-21+1) + (-1^2+ 1^2) * 2^(-2*21) )   n = 21   d_n = -1+1i 
assign X[4'b0111] [21] = 146'h 0000000000000000300000000000000000000;  // -0.0000002384185791 = 0.5 * ln( 1 + -1 * 2^(-22+1) + (-1^2+ 1^2) * 2^(-2*22) )   n = 22   d_n = -1+1i 
assign X[4'b0111] [22] = 146'h 00000000000000000C0000000000000000000;  // -0.0000001192092896 = 0.5 * ln( 1 + -1 * 2^(-23+1) + (-1^2+ 1^2) * 2^(-2*23) )   n = 23   d_n = -1+1i 
assign X[4'b0111] [23] = 146'h 0000000000000000030000000000000000000;  // -0.0000000596046448 = 0.5 * ln( 1 + -1 * 2^(-24+1) + (-1^2+ 1^2) * 2^(-2*24) )   n = 24   d_n = -1+1i 
assign X[4'b0111] [24] = 146'h 000000000000000000C000000000000000000;  // -0.0000000298023224 = 0.5 * ln( 1 + -1 * 2^(-25+1) + (-1^2+ 1^2) * 2^(-2*25) )   n = 25   d_n = -1+1i 
assign X[4'b0111] [25] = 146'h 0000000000000000003000000000000000000;  // -0.0000000149011612 = 0.5 * ln( 1 + -1 * 2^(-26+1) + (-1^2+ 1^2) * 2^(-2*26) )   n = 26   d_n = -1+1i 
assign X[4'b0111] [26] = 146'h 0000000000000000000C00000000000000000;  // -0.0000000074505806 = 0.5 * ln( 1 + -1 * 2^(-27+1) + (-1^2+ 1^2) * 2^(-2*27) )   n = 27   d_n = -1+1i 
assign X[4'b0111] [27] = 146'h 0000000000000000000300000000000000000;  // -0.0000000037252903 = 0.5 * ln( 1 + -1 * 2^(-28+1) + (-1^2+ 1^2) * 2^(-2*28) )   n = 28   d_n = -1+1i 
assign X[4'b0111] [28] = 146'h 00000000000000000000C0000000000000000;  // -0.0000000018626452 = 0.5 * ln( 1 + -1 * 2^(-29+1) + (-1^2+ 1^2) * 2^(-2*29) )   n = 29   d_n = -1+1i 
assign X[4'b0111] [29] = 146'h 0000000000000000000030000000000000000;  // -0.0000000009313226 = 0.5 * ln( 1 + -1 * 2^(-30+1) + (-1^2+ 1^2) * 2^(-2*30) )   n = 30   d_n = -1+1i 
assign X[4'b0111] [30] = 146'h 000000000000000000000C000000000000000;  // -0.0000000004656613 = 0.5 * ln( 1 + -1 * 2^(-31+1) + (-1^2+ 1^2) * 2^(-2*31) )   n = 31   d_n = -1+1i 
assign X[4'b0111] [31] = 146'h 0000000000000000000003000000000000000;  // -0.0000000002328306 = 0.5 * ln( 1 + -1 * 2^(-32+1) + (-1^2+ 1^2) * 2^(-2*32) )   n = 32   d_n = -1+1i 
assign X[4'b0111] [32] = 146'h 0000000000000000000000C00000000000000;  // -0.0000000001164153 = 0.5 * ln( 1 + -1 * 2^(-33+1) + (-1^2+ 1^2) * 2^(-2*33) )   n = 33   d_n = -1+1i 
assign X[4'b0111] [33] = 146'h 0000000000000000000000300000000000000;  // -0.0000000000582077 = 0.5 * ln( 1 + -1 * 2^(-34+1) + (-1^2+ 1^2) * 2^(-2*34) )   n = 34   d_n = -1+1i 
assign X[4'b0111] [34] = 146'h 00000000000000000000000C0000000000000;  // -0.0000000000291038 = 0.5 * ln( 1 + -1 * 2^(-35+1) + (-1^2+ 1^2) * 2^(-2*35) )   n = 35   d_n = -1+1i 
assign X[4'b0111] [35] = 146'h 0000000000000000000000030000000000000;  // -0.0000000000145519 = 0.5 * ln( 1 + -1 * 2^(-36+1) + (-1^2+ 1^2) * 2^(-2*36) )   n = 36   d_n = -1+1i 
assign X[4'b0111] [36] = 146'h 000000000000000000000000C000000000000;  // -0.0000000000072760 = 0.5 * ln( 1 + -1 * 2^(-37+1) + (-1^2+ 1^2) * 2^(-2*37) )   n = 37   d_n = -1+1i 
assign X[4'b0111] [37] = 146'h 0000000000000000000000003000000000000;  // -0.0000000000036380 = 0.5 * ln( 1 + -1 * 2^(-38+1) + (-1^2+ 1^2) * 2^(-2*38) )   n = 38   d_n = -1+1i 
assign X[4'b0111] [38] = 146'h 0000000000000000000000000C00000000000;  // -0.0000000000018190 = 0.5 * ln( 1 + -1 * 2^(-39+1) + (-1^2+ 1^2) * 2^(-2*39) )   n = 39   d_n = -1+1i 
assign X[4'b0111] [39] = 146'h 0000000000000000000000000300000000000;  // -0.0000000000009095 = 0.5 * ln( 1 + -1 * 2^(-40+1) + (-1^2+ 1^2) * 2^(-2*40) )   n = 40   d_n = -1+1i 
assign X[4'b0111] [40] = 146'h 00000000000000000000000000C0000000000;  // -0.0000000000004547 = 0.5 * ln( 1 + -1 * 2^(-41+1) + (-1^2+ 1^2) * 2^(-2*41) )   n = 41   d_n = -1+1i 
assign X[4'b0111] [41] = 146'h 0000000000000000000000000030000000000;  // -0.0000000000002274 = 0.5 * ln( 1 + -1 * 2^(-42+1) + (-1^2+ 1^2) * 2^(-2*42) )   n = 42   d_n = -1+1i 
assign X[4'b0111] [42] = 146'h 000000000000000000000000000C000000000;  // -0.0000000000001137 = 0.5 * ln( 1 + -1 * 2^(-43+1) + (-1^2+ 1^2) * 2^(-2*43) )   n = 43   d_n = -1+1i 
assign X[4'b0111] [43] = 146'h 0000000000000000000000000003000000000;  // -0.0000000000000568 = 0.5 * ln( 1 + -1 * 2^(-44+1) + (-1^2+ 1^2) * 2^(-2*44) )   n = 44   d_n = -1+1i 
assign X[4'b0111] [44] = 146'h 0000000000000000000000000000C00000000;  // -0.0000000000000284 = 0.5 * ln( 1 + -1 * 2^(-45+1) + (-1^2+ 1^2) * 2^(-2*45) )   n = 45   d_n = -1+1i 
assign X[4'b0111] [45] = 146'h 0000000000000000000000000000300000000;  // -0.0000000000000142 = 0.5 * ln( 1 + -1 * 2^(-46+1) + (-1^2+ 1^2) * 2^(-2*46) )   n = 46   d_n = -1+1i 
assign X[4'b0111] [46] = 146'h 00000000000000000000000000000C0000000;  // -0.0000000000000071 = 0.5 * ln( 1 + -1 * 2^(-47+1) + (-1^2+ 1^2) * 2^(-2*47) )   n = 47   d_n = -1+1i 
assign X[4'b0111] [47] = 146'h 0000000000000000000000000000030000000;  // -0.0000000000000036 = 0.5 * ln( 1 + -1 * 2^(-48+1) + (-1^2+ 1^2) * 2^(-2*48) )   n = 48   d_n = -1+1i 
assign X[4'b0111] [48] = 146'h 000000000000000000000000000000C000000;  // -0.0000000000000018 = 0.5 * ln( 1 + -1 * 2^(-49+1) + (-1^2+ 1^2) * 2^(-2*49) )   n = 49   d_n = -1+1i 
assign X[4'b0111] [49] = 146'h 0000000000000000000000000000003000000;  // -0.0000000000000009 = 0.5 * ln( 1 + -1 * 2^(-50+1) + (-1^2+ 1^2) * 2^(-2*50) )   n = 50   d_n = -1+1i 
assign X[4'b0111] [50] = 146'h 0000000000000000000000000000000C00000;  // -0.0000000000000004 = 0.5 * ln( 1 + -1 * 2^(-51+1) + (-1^2+ 1^2) * 2^(-2*51) )   n = 51   d_n = -1+1i 
assign X[4'b0111] [51] = 146'h 0000000000000000000000000000000300000;  // -0.0000000000000002 = 0.5 * ln( 1 + -1 * 2^(-52+1) + (-1^2+ 1^2) * 2^(-2*52) )   n = 52   d_n = -1+1i 
assign X[4'b0111] [52] = 146'h 00000000000000000000000000000000C0000;  // -0.0000000000000001 = 0.5 * ln( 1 + -1 * 2^(-53+1) + (-1^2+ 1^2) * 2^(-2*53) )   n = 53   d_n = -1+1i 
assign X[4'b0111] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-54+1) + (-1^2+ 1^2) * 2^(-2*54) )   n = 54   d_n = -1+1i 
assign X[4'b0111] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-55+1) + (-1^2+ 1^2) * 2^(-2*55) )   n = 55   d_n = -1+1i 
assign X[4'b0111] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-56+1) + (-1^2+ 1^2) * 2^(-2*56) )   n = 56   d_n = -1+1i 
assign X[4'b0111] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-57+1) + (-1^2+ 1^2) * 2^(-2*57) )   n = 57   d_n = -1+1i 
assign X[4'b0111] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-58+1) + (-1^2+ 1^2) * 2^(-2*58) )   n = 58   d_n = -1+1i 
assign X[4'b0111] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-59+1) + (-1^2+ 1^2) * 2^(-2*59) )   n = 59   d_n = -1+1i 
assign X[4'b0111] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-60+1) + (-1^2+ 1^2) * 2^(-2*60) )   n = 60   d_n = -1+1i 
assign X[4'b0111] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-61+1) + (-1^2+ 1^2) * 2^(-2*61) )   n = 61   d_n = -1+1i 
assign X[4'b0111] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-62+1) + (-1^2+ 1^2) * 2^(-2*62) )   n = 62   d_n = -1+1i 
assign X[4'b0111] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-63+1) + (-1^2+ 1^2) * 2^(-2*63) )   n = 63   d_n = -1+1i 
assign X[4'b0111] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-64+1) + (-1^2+ 1^2) * 2^(-2*64) )   n = 64   d_n = -1+1i 
assign X[4'b1000] [00] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-1+1) + ( 0^2+ 0^2) * 2^(-2*1) )   n =  1   d_n = 0 
assign X[4'b1000] [01] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-2+1) + ( 0^2+ 0^2) * 2^(-2*2) )   n =  2   d_n = 0 
assign X[4'b1000] [02] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-3+1) + ( 0^2+ 0^2) * 2^(-2*3) )   n =  3   d_n = 0 
assign X[4'b1000] [03] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-4+1) + ( 0^2+ 0^2) * 2^(-2*4) )   n =  4   d_n = 0 
assign X[4'b1000] [04] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-5+1) + ( 0^2+ 0^2) * 2^(-2*5) )   n =  5   d_n = 0 
assign X[4'b1000] [05] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-6+1) + ( 0^2+ 0^2) * 2^(-2*6) )   n =  6   d_n = 0 
assign X[4'b1000] [06] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-7+1) + ( 0^2+ 0^2) * 2^(-2*7) )   n =  7   d_n = 0 
assign X[4'b1000] [07] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-8+1) + ( 0^2+ 0^2) * 2^(-2*8) )   n =  8   d_n = 0 
assign X[4'b1000] [08] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-9+1) + ( 0^2+ 0^2) * 2^(-2*9) )   n =  9   d_n = 0 
assign X[4'b1000] [09] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = 0 
assign X[4'b1000] [10] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = 0 
assign X[4'b1000] [11] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = 0 
assign X[4'b1000] [12] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = 0 
assign X[4'b1000] [13] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = 0 
assign X[4'b1000] [14] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = 0 
assign X[4'b1000] [15] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = 0 
assign X[4'b1000] [16] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = 0 
assign X[4'b1000] [17] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = 0 
assign X[4'b1000] [18] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = 0 
assign X[4'b1000] [19] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = 0 
assign X[4'b1000] [20] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = 0 
assign X[4'b1000] [21] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = 0 
assign X[4'b1000] [22] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = 0 
assign X[4'b1000] [23] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = 0 
assign X[4'b1000] [24] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = 0 
assign X[4'b1000] [25] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = 0 
assign X[4'b1000] [26] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = 0 
assign X[4'b1000] [27] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = 0 
assign X[4'b1000] [28] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = 0 
assign X[4'b1000] [29] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = 0 
assign X[4'b1000] [30] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = 0 
assign X[4'b1000] [31] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = 0 
assign X[4'b1000] [32] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = 0 
assign X[4'b1000] [33] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = 0 
assign X[4'b1000] [34] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = 0 
assign X[4'b1000] [35] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = 0 
assign X[4'b1000] [36] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = 0 
assign X[4'b1000] [37] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = 0 
assign X[4'b1000] [38] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = 0 
assign X[4'b1000] [39] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = 0 
assign X[4'b1000] [40] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = 0 
assign X[4'b1000] [41] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = 0 
assign X[4'b1000] [42] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = 0 
assign X[4'b1000] [43] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = 0 
assign X[4'b1000] [44] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = 0 
assign X[4'b1000] [45] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = 0 
assign X[4'b1000] [46] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = 0 
assign X[4'b1000] [47] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = 0 
assign X[4'b1000] [48] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = 0 
assign X[4'b1000] [49] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = 0 
assign X[4'b1000] [50] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = 0 
assign X[4'b1000] [51] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = 0 
assign X[4'b1000] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = 0 
assign X[4'b1000] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = 0 
assign X[4'b1000] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = 0 
assign X[4'b1000] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = 0 
assign X[4'b1000] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = 0 
assign X[4'b1000] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = 0 
assign X[4'b1000] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = 0 
assign X[4'b1000] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = 0 
assign X[4'b1000] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = 0 
assign X[4'b1000] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = 0 
assign X[4'b1000] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = 0 
assign X[4'b1000] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = 0 
assign X[4'b1001] [00] = 146'h 0000004C40313041003400000000000000000;  // +0.4054651081081644 = 0.5 * ln( 1 +  1 * 2^(-1+1) + ( 1^2+ 0^2) * 2^(-2*1) )   n =  1   d_n = 1 
assign X[4'b1001] [01] = 146'h 00000010C104000300C100000000000000000;  // +0.2231435513142098 = 0.5 * ln( 1 +  1 * 2^(-2+1) + ( 1^2+ 0^2) * 2^(-2*2) )   n =  2   d_n = 1 
assign X[4'b1001] [02] = 146'h 000000040C04430040C300000000000000000;  // +0.1177830356563835 = 0.5 * ln( 1 +  1 * 2^(-3+1) + ( 1^2+ 0^2) * 2^(-2*3) )   n =  3   d_n = 1 
assign X[4'b1001] [03] = 146'h 0000000100C01104C04C00000000000000000;  // +0.0606246218164348 = 0.5 * ln( 1 +  1 * 2^(-4+1) + ( 1^2+ 0^2) * 2^(-2*4) )   n =  4   d_n = 1 
assign X[4'b1001] [04] = 146'h 00000000400C0044433010000000000000000;  // +0.0307716586667537 = 0.5 * ln( 1 +  1 * 2^(-5+1) + ( 1^2+ 0^2) * 2^(-2*5) )   n =  5   d_n = 1 
assign X[4'b1001] [05] = 146'h 000000001000C0011104CC000000000000000;  // +0.0155041865359653 = 0.5 * ln( 1 +  1 * 2^(-6+1) + ( 1^2+ 0^2) * 2^(-2*6) )   n =  6   d_n = 1 
assign X[4'b1001] [06] = 146'h 0000000004000C00044443400000000000000;  // +0.0077821404420549 = 0.5 * ln( 1 +  1 * 2^(-7+1) + ( 1^2+ 0^2) * 2^(-2*7) )   n =  7   d_n = 1 
assign X[4'b1001] [07] = 146'h 00000000010000C0001111000000000000000;  // +0.0038986404156573 = 0.5 * ln( 1 +  1 * 2^(-8+1) + ( 1^2+ 0^2) * 2^(-2*8) )   n =  8   d_n = 1 
assign X[4'b1001] [08] = 146'h 000000000040000C000044440000000000000;  // +0.0019512201312617 = 0.5 * ln( 1 +  1 * 2^(-9+1) + ( 1^2+ 0^2) * 2^(-2*9) )   n =  9   d_n = 1 
assign X[4'b1001] [09] = 146'h 0000000000100000C00001110000000000000;  // +0.0009760859730555 = 0.5 * ln( 1 +  1 * 2^(-10+1) + ( 1^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = 1 
assign X[4'b1001] [10] = 146'h 00000000000400000C0000044000000000000;  // +0.0004881620795014 = 0.5 * ln( 1 +  1 * 2^(-11+1) + ( 1^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = 1 
assign X[4'b1001] [11] = 146'h 000000000001000000C000001000000000000;  // +0.0002441108275274 = 0.5 * ln( 1 +  1 * 2^(-12+1) + ( 1^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = 1 
assign X[4'b1001] [12] = 146'h 0000000000004000000C00000000000000000;  // +0.0001220628625257 = 0.5 * ln( 1 +  1 * 2^(-13+1) + ( 1^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = 1 
assign X[4'b1001] [13] = 146'h 00000000000010000000C0000000000000000;  // +0.0000610332936806 = 0.5 * ln( 1 +  1 * 2^(-14+1) + ( 1^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = 1 
assign X[4'b1001] [14] = 146'h 000000000000040000000C000000000000000;  // +0.0000305171124732 = 0.5 * ln( 1 +  1 * 2^(-15+1) + ( 1^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = 1 
assign X[4'b1001] [15] = 146'h 0000000000000100000000C00000000000000;  // +0.0000152586726484 = 0.5 * ln( 1 +  1 * 2^(-16+1) + ( 1^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = 1 
assign X[4'b1001] [16] = 146'h 00000000000000400000000C0000000000000;  // +0.0000076293654276 = 0.5 * ln( 1 +  1 * 2^(-17+1) + ( 1^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = 1 
assign X[4'b1001] [17] = 146'h 000000000000001000000000C000000000000;  // +0.0000038146899897 = 0.5 * ln( 1 +  1 * 2^(-18+1) + ( 1^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = 1 
assign X[4'b1001] [18] = 146'h 0000000000000004000000000C00000000000;  // +0.0000019073468138 = 0.5 * ln( 1 +  1 * 2^(-19+1) + ( 1^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = 1 
assign X[4'b1001] [19] = 146'h 00000000000000010000000000C0000000000;  // +0.0000009536738617 = 0.5 * ln( 1 +  1 * 2^(-20+1) + ( 1^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = 1 
assign X[4'b1001] [20] = 146'h 000000000000000040000000000C000000000;  // +0.0000004768370445 = 0.5 * ln( 1 +  1 * 2^(-21+1) + ( 1^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = 1 
assign X[4'b1001] [21] = 146'h 0000000000000000100000000000C00000000;  // +0.0000002384185507 = 0.5 * ln( 1 +  1 * 2^(-22+1) + ( 1^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = 1 
assign X[4'b1001] [22] = 146'h 00000000000000000400000000000C0000000;  // +0.0000001192092824 = 0.5 * ln( 1 +  1 * 2^(-23+1) + ( 1^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = 1 
assign X[4'b1001] [23] = 146'h 000000000000000001000000000000C000000;  // +0.0000000596046430 = 0.5 * ln( 1 +  1 * 2^(-24+1) + ( 1^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = 1 
assign X[4'b1001] [24] = 146'h 0000000000000000004000000000000C00000;  // +0.0000000298023219 = 0.5 * ln( 1 +  1 * 2^(-25+1) + ( 1^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = 1 
assign X[4'b1001] [25] = 146'h 0000000000000000001000000000000100000;  // +0.0000000149011611 = 0.5 * ln( 1 +  1 * 2^(-26+1) + ( 1^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = 1 
assign X[4'b1001] [26] = 146'h 0000000000000000000400000000000000000;  // +0.0000000074505806 = 0.5 * ln( 1 +  1 * 2^(-27+1) + ( 1^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = 1 
assign X[4'b1001] [27] = 146'h 0000000000000000000100000000000000000;  // +0.0000000037252903 = 0.5 * ln( 1 +  1 * 2^(-28+1) + ( 1^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = 1 
assign X[4'b1001] [28] = 146'h 0000000000000000000040000000000000000;  // +0.0000000018626451 = 0.5 * ln( 1 +  1 * 2^(-29+1) + ( 1^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = 1 
assign X[4'b1001] [29] = 146'h 0000000000000000000010000000000000000;  // +0.0000000009313226 = 0.5 * ln( 1 +  1 * 2^(-30+1) + ( 1^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = 1 
assign X[4'b1001] [30] = 146'h 0000000000000000000004000000000000000;  // +0.0000000004656613 = 0.5 * ln( 1 +  1 * 2^(-31+1) + ( 1^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = 1 
assign X[4'b1001] [31] = 146'h 0000000000000000000001000000000000000;  // +0.0000000002328306 = 0.5 * ln( 1 +  1 * 2^(-32+1) + ( 1^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = 1 
assign X[4'b1001] [32] = 146'h 0000000000000000000000400000000000000;  // +0.0000000001164153 = 0.5 * ln( 1 +  1 * 2^(-33+1) + ( 1^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = 1 
assign X[4'b1001] [33] = 146'h 0000000000000000000000100000000000000;  // +0.0000000000582077 = 0.5 * ln( 1 +  1 * 2^(-34+1) + ( 1^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = 1 
assign X[4'b1001] [34] = 146'h 0000000000000000000000040000000000000;  // +0.0000000000291038 = 0.5 * ln( 1 +  1 * 2^(-35+1) + ( 1^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = 1 
assign X[4'b1001] [35] = 146'h 0000000000000000000000010000000000000;  // +0.0000000000145519 = 0.5 * ln( 1 +  1 * 2^(-36+1) + ( 1^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = 1 
assign X[4'b1001] [36] = 146'h 0000000000000000000000004000000000000;  // +0.0000000000072760 = 0.5 * ln( 1 +  1 * 2^(-37+1) + ( 1^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = 1 
assign X[4'b1001] [37] = 146'h 0000000000000000000000001000000000000;  // +0.0000000000036380 = 0.5 * ln( 1 +  1 * 2^(-38+1) + ( 1^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = 1 
assign X[4'b1001] [38] = 146'h 0000000000000000000000000400000000000;  // +0.0000000000018190 = 0.5 * ln( 1 +  1 * 2^(-39+1) + ( 1^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = 1 
assign X[4'b1001] [39] = 146'h 0000000000000000000000000100000000000;  // +0.0000000000009095 = 0.5 * ln( 1 +  1 * 2^(-40+1) + ( 1^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = 1 
assign X[4'b1001] [40] = 146'h 0000000000000000000000000040000000000;  // +0.0000000000004547 = 0.5 * ln( 1 +  1 * 2^(-41+1) + ( 1^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = 1 
assign X[4'b1001] [41] = 146'h 0000000000000000000000000010000000000;  // +0.0000000000002274 = 0.5 * ln( 1 +  1 * 2^(-42+1) + ( 1^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = 1 
assign X[4'b1001] [42] = 146'h 0000000000000000000000000004000000000;  // +0.0000000000001137 = 0.5 * ln( 1 +  1 * 2^(-43+1) + ( 1^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = 1 
assign X[4'b1001] [43] = 146'h 0000000000000000000000000001000000000;  // +0.0000000000000568 = 0.5 * ln( 1 +  1 * 2^(-44+1) + ( 1^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = 1 
assign X[4'b1001] [44] = 146'h 0000000000000000000000000000400000000;  // +0.0000000000000284 = 0.5 * ln( 1 +  1 * 2^(-45+1) + ( 1^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = 1 
assign X[4'b1001] [45] = 146'h 0000000000000000000000000000100000000;  // +0.0000000000000142 = 0.5 * ln( 1 +  1 * 2^(-46+1) + ( 1^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = 1 
assign X[4'b1001] [46] = 146'h 0000000000000000000000000000040000000;  // +0.0000000000000071 = 0.5 * ln( 1 +  1 * 2^(-47+1) + ( 1^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = 1 
assign X[4'b1001] [47] = 146'h 0000000000000000000000000000010000000;  // +0.0000000000000036 = 0.5 * ln( 1 +  1 * 2^(-48+1) + ( 1^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = 1 
assign X[4'b1001] [48] = 146'h 0000000000000000000000000000004000000;  // +0.0000000000000018 = 0.5 * ln( 1 +  1 * 2^(-49+1) + ( 1^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = 1 
assign X[4'b1001] [49] = 146'h 0000000000000000000000000000001000000;  // +0.0000000000000009 = 0.5 * ln( 1 +  1 * 2^(-50+1) + ( 1^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = 1 
assign X[4'b1001] [50] = 146'h 0000000000000000000000000000000400000;  // +0.0000000000000004 = 0.5 * ln( 1 +  1 * 2^(-51+1) + ( 1^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = 1 
assign X[4'b1001] [51] = 146'h 0000000000000000000000000000000100000;  // +0.0000000000000002 = 0.5 * ln( 1 +  1 * 2^(-52+1) + ( 1^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = 1 
assign X[4'b1001] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-53+1) + ( 1^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = 1 
assign X[4'b1001] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-54+1) + ( 1^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = 1 
assign X[4'b1001] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-55+1) + ( 1^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = 1 
assign X[4'b1001] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-56+1) + ( 1^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = 1 
assign X[4'b1001] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-57+1) + ( 1^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = 1 
assign X[4'b1001] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-58+1) + ( 1^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = 1 
assign X[4'b1001] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-59+1) + ( 1^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = 1 
assign X[4'b1001] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-60+1) + ( 1^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = 1 
assign X[4'b1001] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-61+1) + ( 1^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = 1 
assign X[4'b1001] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-62+1) + ( 1^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = 1 
assign X[4'b1001] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-63+1) + ( 1^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = 1 
assign X[4'b1001] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-64+1) + ( 1^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = 1 
assign X[4'b1010] [00] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-1+1) + ( 0^2+ 0^2) * 2^(-2*1) )   n =  1   d_n = -0 
assign X[4'b1010] [01] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-2+1) + ( 0^2+ 0^2) * 2^(-2*2) )   n =  2   d_n = -0 
assign X[4'b1010] [02] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-3+1) + ( 0^2+ 0^2) * 2^(-2*3) )   n =  3   d_n = -0 
assign X[4'b1010] [03] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-4+1) + ( 0^2+ 0^2) * 2^(-2*4) )   n =  4   d_n = -0 
assign X[4'b1010] [04] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-5+1) + ( 0^2+ 0^2) * 2^(-2*5) )   n =  5   d_n = -0 
assign X[4'b1010] [05] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-6+1) + ( 0^2+ 0^2) * 2^(-2*6) )   n =  6   d_n = -0 
assign X[4'b1010] [06] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-7+1) + ( 0^2+ 0^2) * 2^(-2*7) )   n =  7   d_n = -0 
assign X[4'b1010] [07] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-8+1) + ( 0^2+ 0^2) * 2^(-2*8) )   n =  8   d_n = -0 
assign X[4'b1010] [08] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-9+1) + ( 0^2+ 0^2) * 2^(-2*9) )   n =  9   d_n = -0 
assign X[4'b1010] [09] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = -0 
assign X[4'b1010] [10] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = -0 
assign X[4'b1010] [11] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = -0 
assign X[4'b1010] [12] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = -0 
assign X[4'b1010] [13] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = -0 
assign X[4'b1010] [14] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = -0 
assign X[4'b1010] [15] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = -0 
assign X[4'b1010] [16] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = -0 
assign X[4'b1010] [17] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = -0 
assign X[4'b1010] [18] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = -0 
assign X[4'b1010] [19] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = -0 
assign X[4'b1010] [20] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = -0 
assign X[4'b1010] [21] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = -0 
assign X[4'b1010] [22] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = -0 
assign X[4'b1010] [23] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = -0 
assign X[4'b1010] [24] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = -0 
assign X[4'b1010] [25] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = -0 
assign X[4'b1010] [26] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = -0 
assign X[4'b1010] [27] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = -0 
assign X[4'b1010] [28] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = -0 
assign X[4'b1010] [29] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = -0 
assign X[4'b1010] [30] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = -0 
assign X[4'b1010] [31] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = -0 
assign X[4'b1010] [32] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = -0 
assign X[4'b1010] [33] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = -0 
assign X[4'b1010] [34] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = -0 
assign X[4'b1010] [35] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = -0 
assign X[4'b1010] [36] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = -0 
assign X[4'b1010] [37] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = -0 
assign X[4'b1010] [38] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = -0 
assign X[4'b1010] [39] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = -0 
assign X[4'b1010] [40] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = -0 
assign X[4'b1010] [41] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = -0 
assign X[4'b1010] [42] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = -0 
assign X[4'b1010] [43] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = -0 
assign X[4'b1010] [44] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = -0 
assign X[4'b1010] [45] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = -0 
assign X[4'b1010] [46] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = -0 
assign X[4'b1010] [47] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = -0 
assign X[4'b1010] [48] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = -0 
assign X[4'b1010] [49] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = -0 
assign X[4'b1010] [50] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = -0 
assign X[4'b1010] [51] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = -0 
assign X[4'b1010] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = -0 
assign X[4'b1010] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = -0 
assign X[4'b1010] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = -0 
assign X[4'b1010] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = -0 
assign X[4'b1010] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = -0 
assign X[4'b1010] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = -0 
assign X[4'b1010] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = -0 
assign X[4'b1010] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = -0 
assign X[4'b1010] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = -0 
assign X[4'b1010] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = -0 
assign X[4'b1010] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = -0 
assign X[4'b1010] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = -0 
assign X[4'b1011] [00] = 146'h 000003110C410C0C400000000000000000000;  // -0.6931471805599453 = 0.5 * ln( 1 + -1 * 2^(-1+1) + (-1^2+ 0^2) * 2^(-2*1) )   n =  1   d_n = -1 
assign X[4'b1011] [01] = 146'h 00000030CC4CC440C03000000000000000000;  // -0.2876820724517809 = 0.5 * ln( 1 + -1 * 2^(-2+1) + (-1^2+ 0^2) * 2^(-2*2) )   n =  2   d_n = -1 
assign X[4'b1011] [02] = 146'h 0000000C0C31010C130000000000000000000;  // -0.1335313926245226 = 0.5 * ln( 1 + -1 * 2^(-3+1) + (-1^2+ 0^2) * 2^(-2*3) )   n =  3   d_n = -1 
assign X[4'b1011] [03] = 146'h 0000000300C0C44C431040000000000000000;  // -0.0645385211375712 = 0.5 * ln( 1 + -1 * 2^(-4+1) + (-1^2+ 0^2) * 2^(-2*4) )   n =  4   d_n = -1 
assign X[4'b1011] [04] = 146'h 00000000C00C0311011030000000000000000;  // -0.0317486983145803 = 0.5 * ln( 1 + -1 * 2^(-5+1) + (-1^2+ 0^2) * 2^(-2*5) )   n =  5   d_n = -1 
assign X[4'b1011] [05] = 146'h 000000003000C00C444C44000000000000000;  // -0.0157483569681392 = 0.5 * ln( 1 + -1 * 2^(-6+1) + (-1^2+ 0^2) * 2^(-2*6) )   n =  6   d_n = -1 
assign X[4'b1011] [06] = 146'h 000000000C000C00311101000000000000000;  // -0.0078431774610259 = 0.5 * ln( 1 + -1 * 2^(-7+1) + (-1^2+ 0^2) * 2^(-2*7) )   n =  7   d_n = -1 
assign X[4'b1011] [07] = 146'h 00000000030000C000C444400000000000000;  // -0.0039138993211363 = 0.5 * ln( 1 + -1 * 2^(-8+1) + (-1^2+ 0^2) * 2^(-2*8) )   n =  8   d_n = -1 
assign X[4'b1011] [08] = 146'h 0000000000C0000C000311100000000000000;  // -0.0019550348358034 = 0.5 * ln( 1 + -1 * 2^(-9+1) + (-1^2+ 0^2) * 2^(-2*9) )   n =  9   d_n = -1 
assign X[4'b1011] [09] = 146'h 0000000000300000C0000C440000000000000;  // -0.0009770396478266 = 0.5 * ln( 1 + -1 * 2^(-10+1) + (-1^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = -1 
assign X[4'b1011] [10] = 146'h 00000000000C00000C0000310000000000000;  // -0.0004884004981089 = 0.5 * ln( 1 + -1 * 2^(-11+1) + (-1^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = -1 
assign X[4'b1011] [11] = 146'h 000000000003000000C00000C000000000000;  // -0.0002441704321739 = 0.5 * ln( 1 + -1 * 2^(-12+1) + (-1^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = -1 
assign X[4'b1011] [12] = 146'h 000000000000C000000C00000000000000000;  // -0.0001220777636870 = 0.5 * ln( 1 + -1 * 2^(-13+1) + (-1^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = -1 
assign X[4'b1011] [13] = 146'h 00000000000030000000C0000000000000000;  // -0.0000610370189709 = 0.5 * ln( 1 + -1 * 2^(-14+1) + (-1^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = -1 
assign X[4'b1011] [14] = 146'h 0000000000000C0000000C000000000000000;  // -0.0000305180437958 = 0.5 * ln( 1 + -1 * 2^(-15+1) + (-1^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = -1 
assign X[4'b1011] [15] = 146'h 0000000000000300000000C00000000000000;  // -0.0000152589054790 = 0.5 * ln( 1 + -1 * 2^(-16+1) + (-1^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = -1 
assign X[4'b1011] [16] = 146'h 00000000000000C00000000C0000000000000;  // -0.0000076294236352 = 0.5 * ln( 1 + -1 * 2^(-17+1) + (-1^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = -1 
assign X[4'b1011] [17] = 146'h 000000000000003000000000C000000000000;  // -0.0000038147045416 = 0.5 * ln( 1 + -1 * 2^(-18+1) + (-1^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = -1 
assign X[4'b1011] [18] = 146'h 000000000000000C000000000C00000000000;  // -0.0000019073504518 = 0.5 * ln( 1 + -1 * 2^(-19+1) + (-1^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = -1 
assign X[4'b1011] [19] = 146'h 00000000000000030000000000C0000000000;  // -0.0000009536747712 = 0.5 * ln( 1 + -1 * 2^(-20+1) + (-1^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = -1 
assign X[4'b1011] [20] = 146'h 0000000000000000C0000000000C000000000;  // -0.0000004768372719 = 0.5 * ln( 1 + -1 * 2^(-21+1) + (-1^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = -1 
assign X[4'b1011] [21] = 146'h 0000000000000000300000000000C00000000;  // -0.0000002384186075 = 0.5 * ln( 1 + -1 * 2^(-22+1) + (-1^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = -1 
assign X[4'b1011] [22] = 146'h 00000000000000000C00000000000C0000000;  // -0.0000001192092967 = 0.5 * ln( 1 + -1 * 2^(-23+1) + (-1^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = -1 
assign X[4'b1011] [23] = 146'h 000000000000000003000000000000C000000;  // -0.0000000596046466 = 0.5 * ln( 1 + -1 * 2^(-24+1) + (-1^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = -1 
assign X[4'b1011] [24] = 146'h 000000000000000000C000000000001000000;  // -0.0000000298023228 = 0.5 * ln( 1 + -1 * 2^(-25+1) + (-1^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = -1 
assign X[4'b1011] [25] = 146'h 0000000000000000003000000000000000000;  // -0.0000000149011613 = 0.5 * ln( 1 + -1 * 2^(-26+1) + (-1^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = -1 
assign X[4'b1011] [26] = 146'h 0000000000000000000C00000000000000000;  // -0.0000000074505806 = 0.5 * ln( 1 + -1 * 2^(-27+1) + (-1^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = -1 
assign X[4'b1011] [27] = 146'h 0000000000000000000300000000000000000;  // -0.0000000037252903 = 0.5 * ln( 1 + -1 * 2^(-28+1) + (-1^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = -1 
assign X[4'b1011] [28] = 146'h 00000000000000000000C0000000000000000;  // -0.0000000018626452 = 0.5 * ln( 1 + -1 * 2^(-29+1) + (-1^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = -1 
assign X[4'b1011] [29] = 146'h 0000000000000000000030000000000000000;  // -0.0000000009313226 = 0.5 * ln( 1 + -1 * 2^(-30+1) + (-1^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = -1 
assign X[4'b1011] [30] = 146'h 000000000000000000000C000000000000000;  // -0.0000000004656613 = 0.5 * ln( 1 + -1 * 2^(-31+1) + (-1^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = -1 
assign X[4'b1011] [31] = 146'h 0000000000000000000003000000000000000;  // -0.0000000002328306 = 0.5 * ln( 1 + -1 * 2^(-32+1) + (-1^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = -1 
assign X[4'b1011] [32] = 146'h 0000000000000000000000C00000000000000;  // -0.0000000001164153 = 0.5 * ln( 1 + -1 * 2^(-33+1) + (-1^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = -1 
assign X[4'b1011] [33] = 146'h 0000000000000000000000300000000000000;  // -0.0000000000582077 = 0.5 * ln( 1 + -1 * 2^(-34+1) + (-1^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = -1 
assign X[4'b1011] [34] = 146'h 00000000000000000000000C0000000000000;  // -0.0000000000291038 = 0.5 * ln( 1 + -1 * 2^(-35+1) + (-1^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = -1 
assign X[4'b1011] [35] = 146'h 0000000000000000000000030000000000000;  // -0.0000000000145519 = 0.5 * ln( 1 + -1 * 2^(-36+1) + (-1^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = -1 
assign X[4'b1011] [36] = 146'h 000000000000000000000000C000000000000;  // -0.0000000000072760 = 0.5 * ln( 1 + -1 * 2^(-37+1) + (-1^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = -1 
assign X[4'b1011] [37] = 146'h 0000000000000000000000003000000000000;  // -0.0000000000036380 = 0.5 * ln( 1 + -1 * 2^(-38+1) + (-1^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = -1 
assign X[4'b1011] [38] = 146'h 0000000000000000000000000C00000000000;  // -0.0000000000018190 = 0.5 * ln( 1 + -1 * 2^(-39+1) + (-1^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = -1 
assign X[4'b1011] [39] = 146'h 0000000000000000000000000300000000000;  // -0.0000000000009095 = 0.5 * ln( 1 + -1 * 2^(-40+1) + (-1^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = -1 
assign X[4'b1011] [40] = 146'h 00000000000000000000000000C0000000000;  // -0.0000000000004547 = 0.5 * ln( 1 + -1 * 2^(-41+1) + (-1^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = -1 
assign X[4'b1011] [41] = 146'h 0000000000000000000000000030000000000;  // -0.0000000000002274 = 0.5 * ln( 1 + -1 * 2^(-42+1) + (-1^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = -1 
assign X[4'b1011] [42] = 146'h 000000000000000000000000000C000000000;  // -0.0000000000001137 = 0.5 * ln( 1 + -1 * 2^(-43+1) + (-1^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = -1 
assign X[4'b1011] [43] = 146'h 0000000000000000000000000003000000000;  // -0.0000000000000568 = 0.5 * ln( 1 + -1 * 2^(-44+1) + (-1^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = -1 
assign X[4'b1011] [44] = 146'h 0000000000000000000000000000C00000000;  // -0.0000000000000284 = 0.5 * ln( 1 + -1 * 2^(-45+1) + (-1^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = -1 
assign X[4'b1011] [45] = 146'h 0000000000000000000000000000300000000;  // -0.0000000000000142 = 0.5 * ln( 1 + -1 * 2^(-46+1) + (-1^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = -1 
assign X[4'b1011] [46] = 146'h 00000000000000000000000000000C0000000;  // -0.0000000000000071 = 0.5 * ln( 1 + -1 * 2^(-47+1) + (-1^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = -1 
assign X[4'b1011] [47] = 146'h 0000000000000000000000000000030000000;  // -0.0000000000000036 = 0.5 * ln( 1 + -1 * 2^(-48+1) + (-1^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = -1 
assign X[4'b1011] [48] = 146'h 000000000000000000000000000000C000000;  // -0.0000000000000018 = 0.5 * ln( 1 + -1 * 2^(-49+1) + (-1^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = -1 
assign X[4'b1011] [49] = 146'h 0000000000000000000000000000003000000;  // -0.0000000000000009 = 0.5 * ln( 1 + -1 * 2^(-50+1) + (-1^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = -1 
assign X[4'b1011] [50] = 146'h 0000000000000000000000000000000C00000;  // -0.0000000000000004 = 0.5 * ln( 1 + -1 * 2^(-51+1) + (-1^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = -1 
assign X[4'b1011] [51] = 146'h 0000000000000000000000000000000300000;  // -0.0000000000000002 = 0.5 * ln( 1 + -1 * 2^(-52+1) + (-1^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = -1 
assign X[4'b1011] [52] = 146'h 00000000000000000000000000000000C0000;  // -0.0000000000000001 = 0.5 * ln( 1 + -1 * 2^(-53+1) + (-1^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = -1 
assign X[4'b1011] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-54+1) + (-1^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = -1 
assign X[4'b1011] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-55+1) + (-1^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = -1 
assign X[4'b1011] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-56+1) + (-1^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = -1 
assign X[4'b1011] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-57+1) + (-1^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = -1 
assign X[4'b1011] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-58+1) + (-1^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = -1 
assign X[4'b1011] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-59+1) + (-1^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = -1 
assign X[4'b1011] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-60+1) + (-1^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = -1 
assign X[4'b1011] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-61+1) + (-1^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = -1 
assign X[4'b1011] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-62+1) + (-1^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = -1 
assign X[4'b1011] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-63+1) + (-1^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = -1 
assign X[4'b1011] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-64+1) + (-1^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = -1 
assign X[4'b1100] [00] = 146'h 0000000430410000C03040000000000000000;  // +0.1115717756571049 = 0.5 * ln( 1 +  0 * 2^(-1+1) + ( 0^2+-1^2) * 2^(-2*1) )   n =  1   d_n = -0-1i 
assign X[4'b1100] [01] = 146'h 0000000040300441301300000000000000000;  // +0.0303123109082174 = 0.5 * ln( 1 +  0 * 2^(-2+1) + ( 0^2+-1^2) * 2^(-2*2) )   n =  2   d_n = -0-1i 
assign X[4'b1100] [02] = 146'h 0000000004003000444133000000000000000;  // +0.0077520932679826 = 0.5 * ln( 1 +  0 * 2^(-3+1) + ( 0^2+-1^2) * 2^(-2*3) )   n =  3   d_n = -0-1i 
assign X[4'b1100] [03] = 146'h 0000000000400030000444400000000000000;  // +0.0019493202078287 = 0.5 * ln( 1 +  0 * 2^(-4+1) + ( 0^2+-1^2) * 2^(-2*4) )   n =  4   d_n = -0-1i 
assign X[4'b1100] [04] = 146'h 0000000000040000300000444000000000000;  // +0.0004880429865277 = 0.5 * ln( 1 +  0 * 2^(-5+1) + ( 0^2+-1^2) * 2^(-2*5) )   n =  5   d_n = -0-1i 
assign X[4'b1100] [05] = 146'h 0000000000004000003000000400000000000;  // +0.0001220554137636 = 0.5 * ln( 1 +  0 * 2^(-6+1) + ( 0^2+-1^2) * 2^(-2*6) )   n =  6   d_n = -0-1i 
assign X[4'b1100] [06] = 146'h 0000000000000400000030000000000000000;  // +0.0000305166468403 = 0.5 * ln( 1 +  0 * 2^(-7+1) + ( 0^2+-1^2) * 2^(-2*7) )   n =  7   d_n = -0-1i 
assign X[4'b1100] [07] = 146'h 0000000000000040000000300000000000000;  // +0.0000076293363242 = 0.5 * ln( 1 +  0 * 2^(-8+1) + ( 0^2+-1^2) * 2^(-2*8) )   n =  8   d_n = -0-1i 
assign X[4'b1100] [08] = 146'h 0000000000000004000000003000000000000;  // +0.0000019073449948 = 0.5 * ln( 1 +  0 * 2^(-9+1) + ( 0^2+-1^2) * 2^(-2*9) )   n =  9   d_n = -0-1i 
assign X[4'b1100] [09] = 146'h 0000000000000000400000000030000000000;  // +0.0000004768369308 = 0.5 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+-1^2) * 2^(-2*10) )   n = 10   d_n = -0-1i 
assign X[4'b1100] [10] = 146'h 0000000000000000040000000000300000000;  // +0.0000001192092753 = 0.5 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+-1^2) * 2^(-2*11) )   n = 11   d_n = -0-1i 
assign X[4'b1100] [11] = 146'h 0000000000000000004000000000003000000;  // +0.0000000298023215 = 0.5 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+-1^2) * 2^(-2*12) )   n = 12   d_n = -0-1i 
assign X[4'b1100] [12] = 146'h 0000000000000000000400000000000000000;  // +0.0000000074505806 = 0.5 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+-1^2) * 2^(-2*13) )   n = 13   d_n = -0-1i 
assign X[4'b1100] [13] = 146'h 0000000000000000000040000000000000000;  // +0.0000000018626451 = 0.5 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+-1^2) * 2^(-2*14) )   n = 14   d_n = -0-1i 
assign X[4'b1100] [14] = 146'h 0000000000000000000004000000000000000;  // +0.0000000004656613 = 0.5 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+-1^2) * 2^(-2*15) )   n = 15   d_n = -0-1i 
assign X[4'b1100] [15] = 146'h 0000000000000000000000400000000000000;  // +0.0000000001164153 = 0.5 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+-1^2) * 2^(-2*16) )   n = 16   d_n = -0-1i 
assign X[4'b1100] [16] = 146'h 0000000000000000000000040000000000000;  // +0.0000000000291038 = 0.5 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+-1^2) * 2^(-2*17) )   n = 17   d_n = -0-1i 
assign X[4'b1100] [17] = 146'h 0000000000000000000000004000000000000;  // +0.0000000000072760 = 0.5 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+-1^2) * 2^(-2*18) )   n = 18   d_n = -0-1i 
assign X[4'b1100] [18] = 146'h 0000000000000000000000000400000000000;  // +0.0000000000018190 = 0.5 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+-1^2) * 2^(-2*19) )   n = 19   d_n = -0-1i 
assign X[4'b1100] [19] = 146'h 0000000000000000000000000040000000000;  // +0.0000000000004547 = 0.5 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+-1^2) * 2^(-2*20) )   n = 20   d_n = -0-1i 
assign X[4'b1100] [20] = 146'h 0000000000000000000000000004000000000;  // +0.0000000000001137 = 0.5 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+-1^2) * 2^(-2*21) )   n = 21   d_n = -0-1i 
assign X[4'b1100] [21] = 146'h 0000000000000000000000000000400000000;  // +0.0000000000000284 = 0.5 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+-1^2) * 2^(-2*22) )   n = 22   d_n = -0-1i 
assign X[4'b1100] [22] = 146'h 0000000000000000000000000000040000000;  // +0.0000000000000071 = 0.5 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+-1^2) * 2^(-2*23) )   n = 23   d_n = -0-1i 
assign X[4'b1100] [23] = 146'h 0000000000000000000000000000004000000;  // +0.0000000000000018 = 0.5 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+-1^2) * 2^(-2*24) )   n = 24   d_n = -0-1i 
assign X[4'b1100] [24] = 146'h 0000000000000000000000000000000400000;  // +0.0000000000000004 = 0.5 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+-1^2) * 2^(-2*25) )   n = 25   d_n = -0-1i 
assign X[4'b1100] [25] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+-1^2) * 2^(-2*26) )   n = 26   d_n = -0-1i 
assign X[4'b1100] [26] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+-1^2) * 2^(-2*27) )   n = 27   d_n = -0-1i 
assign X[4'b1100] [27] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+-1^2) * 2^(-2*28) )   n = 28   d_n = -0-1i 
assign X[4'b1100] [28] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+-1^2) * 2^(-2*29) )   n = 29   d_n = -0-1i 
assign X[4'b1100] [29] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+-1^2) * 2^(-2*30) )   n = 30   d_n = -0-1i 
assign X[4'b1100] [30] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+-1^2) * 2^(-2*31) )   n = 31   d_n = -0-1i 
assign X[4'b1100] [31] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+-1^2) * 2^(-2*32) )   n = 32   d_n = -0-1i 
assign X[4'b1100] [32] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+-1^2) * 2^(-2*33) )   n = 33   d_n = -0-1i 
assign X[4'b1100] [33] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+-1^2) * 2^(-2*34) )   n = 34   d_n = -0-1i 
assign X[4'b1100] [34] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+-1^2) * 2^(-2*35) )   n = 35   d_n = -0-1i 
assign X[4'b1100] [35] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+-1^2) * 2^(-2*36) )   n = 36   d_n = -0-1i 
assign X[4'b1100] [36] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+-1^2) * 2^(-2*37) )   n = 37   d_n = -0-1i 
assign X[4'b1100] [37] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+-1^2) * 2^(-2*38) )   n = 38   d_n = -0-1i 
assign X[4'b1100] [38] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+-1^2) * 2^(-2*39) )   n = 39   d_n = -0-1i 
assign X[4'b1100] [39] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+-1^2) * 2^(-2*40) )   n = 40   d_n = -0-1i 
assign X[4'b1100] [40] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+-1^2) * 2^(-2*41) )   n = 41   d_n = -0-1i 
assign X[4'b1100] [41] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+-1^2) * 2^(-2*42) )   n = 42   d_n = -0-1i 
assign X[4'b1100] [42] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+-1^2) * 2^(-2*43) )   n = 43   d_n = -0-1i 
assign X[4'b1100] [43] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+-1^2) * 2^(-2*44) )   n = 44   d_n = -0-1i 
assign X[4'b1100] [44] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+-1^2) * 2^(-2*45) )   n = 45   d_n = -0-1i 
assign X[4'b1100] [45] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+-1^2) * 2^(-2*46) )   n = 46   d_n = -0-1i 
assign X[4'b1100] [46] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+-1^2) * 2^(-2*47) )   n = 47   d_n = -0-1i 
assign X[4'b1100] [47] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+-1^2) * 2^(-2*48) )   n = 48   d_n = -0-1i 
assign X[4'b1100] [48] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+-1^2) * 2^(-2*49) )   n = 49   d_n = -0-1i 
assign X[4'b1100] [49] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+-1^2) * 2^(-2*50) )   n = 50   d_n = -0-1i 
assign X[4'b1100] [50] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+-1^2) * 2^(-2*51) )   n = 51   d_n = -0-1i 
assign X[4'b1100] [51] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+-1^2) * 2^(-2*52) )   n = 52   d_n = -0-1i 
assign X[4'b1100] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+-1^2) * 2^(-2*53) )   n = 53   d_n = -0-1i 
assign X[4'b1100] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+-1^2) * 2^(-2*54) )   n = 54   d_n = -0-1i 
assign X[4'b1100] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+-1^2) * 2^(-2*55) )   n = 55   d_n = -0-1i 
assign X[4'b1100] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+-1^2) * 2^(-2*56) )   n = 56   d_n = -0-1i 
assign X[4'b1100] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+-1^2) * 2^(-2*57) )   n = 57   d_n = -0-1i 
assign X[4'b1100] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+-1^2) * 2^(-2*58) )   n = 58   d_n = -0-1i 
assign X[4'b1100] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+-1^2) * 2^(-2*59) )   n = 59   d_n = -0-1i 
assign X[4'b1100] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+-1^2) * 2^(-2*60) )   n = 60   d_n = -0-1i 
assign X[4'b1100] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+-1^2) * 2^(-2*61) )   n = 61   d_n = -0-1i 
assign X[4'b1100] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+-1^2) * 2^(-2*62) )   n = 62   d_n = -0-1i 
assign X[4'b1100] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+-1^2) * 2^(-2*63) )   n = 63   d_n = -0-1i 
assign X[4'b1100] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+-1^2) * 2^(-2*64) )   n = 64   d_n = -0-1i 
assign X[4'b1101] [00] = 146'h 0000004311104100103000000000000000000;  // +0.4581453659370776 = 0.5 * ln( 1 +  1 * 2^(-1+1) + ( 1^2+-1^2) * 2^(-2*1) )   n =  1   d_n = 1-1i 
assign X[4'b1101] [01] = 146'h 000000100C041104033000000000000000000;  // +0.2427539078908503 = 0.5 * ln( 1 +  1 * 2^(-2+1) + ( 1^2+-1^2) * 2^(-2*2) )   n =  2   d_n = 1-1i 
assign X[4'b1101] [02] = 146'h 000000040030C104C04300000000000000000;  // +0.1239180819522907 = 0.5 * ln( 1 +  1 * 2^(-3+1) + ( 1^2+-1^2) * 2^(-2*3) )   n =  3   d_n = 1-1i 
assign X[4'b1101] [03] = 146'h 000000010000CC104044C0000000000000000;  // +0.0623517392504787 = 0.5 * ln( 1 +  1 * 2^(-4+1) + ( 1^2+-1^2) * 2^(-2*4) )   n =  4   d_n = 1-1i 
assign X[4'b1101] [04] = 146'h 0000000040000330C41010000000000000000;  // +0.0312305848118681 = 0.5 * ln( 1 +  1 * 2^(-5+1) + ( 1^2+-1^2) * 2^(-2*5) )   n =  5   d_n = 1-1i 
assign X[4'b1101] [05] = 146'h 000000001000000CCC1104000000000000000;  // +0.0156225157283291 = 0.5 * ln( 1 +  1 * 2^(-6+1) + ( 1^2+-1^2) * 2^(-2*6) )   n =  6   d_n = 1-1i 
assign X[4'b1101] [06] = 146'h 00000000040000003330C4400000000000000;  // +0.0078121858105703 = 0.5 * ln( 1 +  1 * 2^(-7+1) + ( 1^2+-1^2) * 2^(-2*7) )   n =  7   d_n = 1-1i 
assign X[4'b1101] [07] = 146'h 000000000100000000CCCC100000000000000;  // +0.0039062104956732 = 0.5 * ln( 1 +  1 * 2^(-8+1) + ( 1^2+-1^2) * 2^(-2*8) )   n =  8   d_n = 1-1i 
assign X[4'b1101] [08] = 146'h 0000000000400000000333300000000000000;  // +0.0019531200474755 = 0.5 * ln( 1 +  1 * 2^(-9+1) + ( 1^2+-1^2) * 2^(-2*9) )   n =  9   d_n = 1-1i 
assign X[4'b1101] [09] = 146'h 000000000010000000000CCD0000000000000;  // +0.0009765618800270 = 0.5 * ln( 1 +  1 * 2^(-10+1) + ( 1^2+-1^2) * 2^(-2*10) )   n = 10   d_n = 1-1i 
assign X[4'b1101] [10] = 146'h 0000000000040000000000334000000000000;  // +0.0004882811724466 = 0.5 * ln( 1 +  1 * 2^(-11+1) + ( 1^2+-1^2) * 2^(-2*11) )   n = 11   d_n = 1-1i 
assign X[4'b1101] [11] = 146'h 000000000001000000000000D000000000000;  // +0.0002441406153023 = 0.5 * ln( 1 +  1 * 2^(-12+1) + ( 1^2+-1^2) * 2^(-2*12) )   n = 12   d_n = 1-1i 
assign X[4'b1101] [12] = 146'h 0000000000004000000000000400000000000;  // +0.0001220703112875 = 0.5 * ln( 1 +  1 * 2^(-13+1) + ( 1^2+-1^2) * 2^(-2*13) )   n = 13   d_n = 1-1i 
assign X[4'b1101] [13] = 146'h 0000000000001000000000000000000000000;  // +0.0000610351560984 = 0.5 * ln( 1 +  1 * 2^(-14+1) + ( 1^2+-1^2) * 2^(-2*14) )   n = 14   d_n = 1-1i 
assign X[4'b1101] [14] = 146'h 0000000000000400000000000000000000000;  // +0.0000305175781061 = 0.5 * ln( 1 +  1 * 2^(-15+1) + ( 1^2+-1^2) * 2^(-2*15) )   n = 15   d_n = 1-1i 
assign X[4'b1101] [15] = 146'h 0000000000000100000000000000000000000;  // +0.0000152587890601 = 0.5 * ln( 1 +  1 * 2^(-16+1) + ( 1^2+-1^2) * 2^(-2*16) )   n = 16   d_n = 1-1i 
assign X[4'b1101] [16] = 146'h 0000000000000040000000000000000000000;  // +0.0000076293945310 = 0.5 * ln( 1 +  1 * 2^(-17+1) + ( 1^2+-1^2) * 2^(-2*17) )   n = 17   d_n = 1-1i 
assign X[4'b1101] [17] = 146'h 0000000000000010000000000000000000000;  // +0.0000038146972656 = 0.5 * ln( 1 +  1 * 2^(-18+1) + ( 1^2+-1^2) * 2^(-2*18) )   n = 18   d_n = 1-1i 
assign X[4'b1101] [18] = 146'h 0000000000000004000000000000000000000;  // +0.0000019073486328 = 0.5 * ln( 1 +  1 * 2^(-19+1) + ( 1^2+-1^2) * 2^(-2*19) )   n = 19   d_n = 1-1i 
assign X[4'b1101] [19] = 146'h 0000000000000001000000000000000000000;  // +0.0000009536743164 = 0.5 * ln( 1 +  1 * 2^(-20+1) + ( 1^2+-1^2) * 2^(-2*20) )   n = 20   d_n = 1-1i 
assign X[4'b1101] [20] = 146'h 0000000000000000400000000000000000000;  // +0.0000004768371582 = 0.5 * ln( 1 +  1 * 2^(-21+1) + ( 1^2+-1^2) * 2^(-2*21) )   n = 21   d_n = 1-1i 
assign X[4'b1101] [21] = 146'h 0000000000000000100000000000000000000;  // +0.0000002384185791 = 0.5 * ln( 1 +  1 * 2^(-22+1) + ( 1^2+-1^2) * 2^(-2*22) )   n = 22   d_n = 1-1i 
assign X[4'b1101] [22] = 146'h 0000000000000000040000000000000000000;  // +0.0000001192092896 = 0.5 * ln( 1 +  1 * 2^(-23+1) + ( 1^2+-1^2) * 2^(-2*23) )   n = 23   d_n = 1-1i 
assign X[4'b1101] [23] = 146'h 0000000000000000010000000000000000000;  // +0.0000000596046448 = 0.5 * ln( 1 +  1 * 2^(-24+1) + ( 1^2+-1^2) * 2^(-2*24) )   n = 24   d_n = 1-1i 
assign X[4'b1101] [24] = 146'h 0000000000000000004000000000000000000;  // +0.0000000298023224 = 0.5 * ln( 1 +  1 * 2^(-25+1) + ( 1^2+-1^2) * 2^(-2*25) )   n = 25   d_n = 1-1i 
assign X[4'b1101] [25] = 146'h 0000000000000000001000000000000100000;  // +0.0000000149011611 = 0.5 * ln( 1 +  1 * 2^(-26+1) + ( 1^2+-1^2) * 2^(-2*26) )   n = 26   d_n = 1-1i 
assign X[4'b1101] [26] = 146'h 0000000000000000000400000000000000000;  // +0.0000000074505806 = 0.5 * ln( 1 +  1 * 2^(-27+1) + ( 1^2+-1^2) * 2^(-2*27) )   n = 27   d_n = 1-1i 
assign X[4'b1101] [27] = 146'h 0000000000000000000100000000000000000;  // +0.0000000037252903 = 0.5 * ln( 1 +  1 * 2^(-28+1) + ( 1^2+-1^2) * 2^(-2*28) )   n = 28   d_n = 1-1i 
assign X[4'b1101] [28] = 146'h 0000000000000000000040000000000000000;  // +0.0000000018626451 = 0.5 * ln( 1 +  1 * 2^(-29+1) + ( 1^2+-1^2) * 2^(-2*29) )   n = 29   d_n = 1-1i 
assign X[4'b1101] [29] = 146'h 0000000000000000000010000000000000000;  // +0.0000000009313226 = 0.5 * ln( 1 +  1 * 2^(-30+1) + ( 1^2+-1^2) * 2^(-2*30) )   n = 30   d_n = 1-1i 
assign X[4'b1101] [30] = 146'h 0000000000000000000004000000000000000;  // +0.0000000004656613 = 0.5 * ln( 1 +  1 * 2^(-31+1) + ( 1^2+-1^2) * 2^(-2*31) )   n = 31   d_n = 1-1i 
assign X[4'b1101] [31] = 146'h 0000000000000000000001000000000000000;  // +0.0000000002328306 = 0.5 * ln( 1 +  1 * 2^(-32+1) + ( 1^2+-1^2) * 2^(-2*32) )   n = 32   d_n = 1-1i 
assign X[4'b1101] [32] = 146'h 0000000000000000000000400000000000000;  // +0.0000000001164153 = 0.5 * ln( 1 +  1 * 2^(-33+1) + ( 1^2+-1^2) * 2^(-2*33) )   n = 33   d_n = 1-1i 
assign X[4'b1101] [33] = 146'h 0000000000000000000000100000000000000;  // +0.0000000000582077 = 0.5 * ln( 1 +  1 * 2^(-34+1) + ( 1^2+-1^2) * 2^(-2*34) )   n = 34   d_n = 1-1i 
assign X[4'b1101] [34] = 146'h 0000000000000000000000040000000000000;  // +0.0000000000291038 = 0.5 * ln( 1 +  1 * 2^(-35+1) + ( 1^2+-1^2) * 2^(-2*35) )   n = 35   d_n = 1-1i 
assign X[4'b1101] [35] = 146'h 0000000000000000000000010000000000000;  // +0.0000000000145519 = 0.5 * ln( 1 +  1 * 2^(-36+1) + ( 1^2+-1^2) * 2^(-2*36) )   n = 36   d_n = 1-1i 
assign X[4'b1101] [36] = 146'h 0000000000000000000000004000000000000;  // +0.0000000000072760 = 0.5 * ln( 1 +  1 * 2^(-37+1) + ( 1^2+-1^2) * 2^(-2*37) )   n = 37   d_n = 1-1i 
assign X[4'b1101] [37] = 146'h 0000000000000000000000001000000000000;  // +0.0000000000036380 = 0.5 * ln( 1 +  1 * 2^(-38+1) + ( 1^2+-1^2) * 2^(-2*38) )   n = 38   d_n = 1-1i 
assign X[4'b1101] [38] = 146'h 0000000000000000000000000400000000000;  // +0.0000000000018190 = 0.5 * ln( 1 +  1 * 2^(-39+1) + ( 1^2+-1^2) * 2^(-2*39) )   n = 39   d_n = 1-1i 
assign X[4'b1101] [39] = 146'h 0000000000000000000000000100000000000;  // +0.0000000000009095 = 0.5 * ln( 1 +  1 * 2^(-40+1) + ( 1^2+-1^2) * 2^(-2*40) )   n = 40   d_n = 1-1i 
assign X[4'b1101] [40] = 146'h 0000000000000000000000000040000000000;  // +0.0000000000004547 = 0.5 * ln( 1 +  1 * 2^(-41+1) + ( 1^2+-1^2) * 2^(-2*41) )   n = 41   d_n = 1-1i 
assign X[4'b1101] [41] = 146'h 0000000000000000000000000010000000000;  // +0.0000000000002274 = 0.5 * ln( 1 +  1 * 2^(-42+1) + ( 1^2+-1^2) * 2^(-2*42) )   n = 42   d_n = 1-1i 
assign X[4'b1101] [42] = 146'h 0000000000000000000000000004000000000;  // +0.0000000000001137 = 0.5 * ln( 1 +  1 * 2^(-43+1) + ( 1^2+-1^2) * 2^(-2*43) )   n = 43   d_n = 1-1i 
assign X[4'b1101] [43] = 146'h 0000000000000000000000000001000000000;  // +0.0000000000000568 = 0.5 * ln( 1 +  1 * 2^(-44+1) + ( 1^2+-1^2) * 2^(-2*44) )   n = 44   d_n = 1-1i 
assign X[4'b1101] [44] = 146'h 0000000000000000000000000000400000000;  // +0.0000000000000284 = 0.5 * ln( 1 +  1 * 2^(-45+1) + ( 1^2+-1^2) * 2^(-2*45) )   n = 45   d_n = 1-1i 
assign X[4'b1101] [45] = 146'h 0000000000000000000000000000100000000;  // +0.0000000000000142 = 0.5 * ln( 1 +  1 * 2^(-46+1) + ( 1^2+-1^2) * 2^(-2*46) )   n = 46   d_n = 1-1i 
assign X[4'b1101] [46] = 146'h 0000000000000000000000000000040000000;  // +0.0000000000000071 = 0.5 * ln( 1 +  1 * 2^(-47+1) + ( 1^2+-1^2) * 2^(-2*47) )   n = 47   d_n = 1-1i 
assign X[4'b1101] [47] = 146'h 0000000000000000000000000000010000000;  // +0.0000000000000036 = 0.5 * ln( 1 +  1 * 2^(-48+1) + ( 1^2+-1^2) * 2^(-2*48) )   n = 48   d_n = 1-1i 
assign X[4'b1101] [48] = 146'h 0000000000000000000000000000004000000;  // +0.0000000000000018 = 0.5 * ln( 1 +  1 * 2^(-49+1) + ( 1^2+-1^2) * 2^(-2*49) )   n = 49   d_n = 1-1i 
assign X[4'b1101] [49] = 146'h 0000000000000000000000000000001000000;  // +0.0000000000000009 = 0.5 * ln( 1 +  1 * 2^(-50+1) + ( 1^2+-1^2) * 2^(-2*50) )   n = 50   d_n = 1-1i 
assign X[4'b1101] [50] = 146'h 0000000000000000000000000000000400000;  // +0.0000000000000004 = 0.5 * ln( 1 +  1 * 2^(-51+1) + ( 1^2+-1^2) * 2^(-2*51) )   n = 51   d_n = 1-1i 
assign X[4'b1101] [51] = 146'h 0000000000000000000000000000000100000;  // +0.0000000000000002 = 0.5 * ln( 1 +  1 * 2^(-52+1) + ( 1^2+-1^2) * 2^(-2*52) )   n = 52   d_n = 1-1i 
assign X[4'b1101] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-53+1) + ( 1^2+-1^2) * 2^(-2*53) )   n = 53   d_n = 1-1i 
assign X[4'b1101] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-54+1) + ( 1^2+-1^2) * 2^(-2*54) )   n = 54   d_n = 1-1i 
assign X[4'b1101] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-55+1) + ( 1^2+-1^2) * 2^(-2*55) )   n = 55   d_n = 1-1i 
assign X[4'b1101] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-56+1) + ( 1^2+-1^2) * 2^(-2*56) )   n = 56   d_n = 1-1i 
assign X[4'b1101] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-57+1) + ( 1^2+-1^2) * 2^(-2*57) )   n = 57   d_n = 1-1i 
assign X[4'b1101] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-58+1) + ( 1^2+-1^2) * 2^(-2*58) )   n = 58   d_n = 1-1i 
assign X[4'b1101] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-59+1) + ( 1^2+-1^2) * 2^(-2*59) )   n = 59   d_n = 1-1i 
assign X[4'b1101] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-60+1) + ( 1^2+-1^2) * 2^(-2*60) )   n = 60   d_n = 1-1i 
assign X[4'b1101] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-61+1) + ( 1^2+-1^2) * 2^(-2*61) )   n = 61   d_n = 1-1i 
assign X[4'b1101] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-62+1) + ( 1^2+-1^2) * 2^(-2*62) )   n = 62   d_n = 1-1i 
assign X[4'b1101] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-63+1) + ( 1^2+-1^2) * 2^(-2*63) )   n = 63   d_n = 1-1i 
assign X[4'b1101] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-64+1) + ( 1^2+-1^2) * 2^(-2*64) )   n = 64   d_n = 1-1i 
assign X[4'b1110] [00] = 146'h 0000000430410000C03040000000000000000;  // +0.1115717756571049 = 0.5 * ln( 1 +  0 * 2^(-1+1) + ( 0^2+-1^2) * 2^(-2*1) )   n =  1   d_n = -0-1i 
assign X[4'b1110] [01] = 146'h 0000000040300441301300000000000000000;  // +0.0303123109082174 = 0.5 * ln( 1 +  0 * 2^(-2+1) + ( 0^2+-1^2) * 2^(-2*2) )   n =  2   d_n = -0-1i 
assign X[4'b1110] [02] = 146'h 0000000004003000444133000000000000000;  // +0.0077520932679826 = 0.5 * ln( 1 +  0 * 2^(-3+1) + ( 0^2+-1^2) * 2^(-2*3) )   n =  3   d_n = -0-1i 
assign X[4'b1110] [03] = 146'h 0000000000400030000444400000000000000;  // +0.0019493202078287 = 0.5 * ln( 1 +  0 * 2^(-4+1) + ( 0^2+-1^2) * 2^(-2*4) )   n =  4   d_n = -0-1i 
assign X[4'b1110] [04] = 146'h 0000000000040000300000444000000000000;  // +0.0004880429865277 = 0.5 * ln( 1 +  0 * 2^(-5+1) + ( 0^2+-1^2) * 2^(-2*5) )   n =  5   d_n = -0-1i 
assign X[4'b1110] [05] = 146'h 0000000000004000003000000400000000000;  // +0.0001220554137636 = 0.5 * ln( 1 +  0 * 2^(-6+1) + ( 0^2+-1^2) * 2^(-2*6) )   n =  6   d_n = -0-1i 
assign X[4'b1110] [06] = 146'h 0000000000000400000030000000000000000;  // +0.0000305166468403 = 0.5 * ln( 1 +  0 * 2^(-7+1) + ( 0^2+-1^2) * 2^(-2*7) )   n =  7   d_n = -0-1i 
assign X[4'b1110] [07] = 146'h 0000000000000040000000300000000000000;  // +0.0000076293363242 = 0.5 * ln( 1 +  0 * 2^(-8+1) + ( 0^2+-1^2) * 2^(-2*8) )   n =  8   d_n = -0-1i 
assign X[4'b1110] [08] = 146'h 0000000000000004000000003000000000000;  // +0.0000019073449948 = 0.5 * ln( 1 +  0 * 2^(-9+1) + ( 0^2+-1^2) * 2^(-2*9) )   n =  9   d_n = -0-1i 
assign X[4'b1110] [09] = 146'h 0000000000000000400000000030000000000;  // +0.0000004768369308 = 0.5 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+-1^2) * 2^(-2*10) )   n = 10   d_n = -0-1i 
assign X[4'b1110] [10] = 146'h 0000000000000000040000000000300000000;  // +0.0000001192092753 = 0.5 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+-1^2) * 2^(-2*11) )   n = 11   d_n = -0-1i 
assign X[4'b1110] [11] = 146'h 0000000000000000004000000000003000000;  // +0.0000000298023215 = 0.5 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+-1^2) * 2^(-2*12) )   n = 12   d_n = -0-1i 
assign X[4'b1110] [12] = 146'h 0000000000000000000400000000000000000;  // +0.0000000074505806 = 0.5 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+-1^2) * 2^(-2*13) )   n = 13   d_n = -0-1i 
assign X[4'b1110] [13] = 146'h 0000000000000000000040000000000000000;  // +0.0000000018626451 = 0.5 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+-1^2) * 2^(-2*14) )   n = 14   d_n = -0-1i 
assign X[4'b1110] [14] = 146'h 0000000000000000000004000000000000000;  // +0.0000000004656613 = 0.5 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+-1^2) * 2^(-2*15) )   n = 15   d_n = -0-1i 
assign X[4'b1110] [15] = 146'h 0000000000000000000000400000000000000;  // +0.0000000001164153 = 0.5 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+-1^2) * 2^(-2*16) )   n = 16   d_n = -0-1i 
assign X[4'b1110] [16] = 146'h 0000000000000000000000040000000000000;  // +0.0000000000291038 = 0.5 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+-1^2) * 2^(-2*17) )   n = 17   d_n = -0-1i 
assign X[4'b1110] [17] = 146'h 0000000000000000000000004000000000000;  // +0.0000000000072760 = 0.5 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+-1^2) * 2^(-2*18) )   n = 18   d_n = -0-1i 
assign X[4'b1110] [18] = 146'h 0000000000000000000000000400000000000;  // +0.0000000000018190 = 0.5 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+-1^2) * 2^(-2*19) )   n = 19   d_n = -0-1i 
assign X[4'b1110] [19] = 146'h 0000000000000000000000000040000000000;  // +0.0000000000004547 = 0.5 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+-1^2) * 2^(-2*20) )   n = 20   d_n = -0-1i 
assign X[4'b1110] [20] = 146'h 0000000000000000000000000004000000000;  // +0.0000000000001137 = 0.5 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+-1^2) * 2^(-2*21) )   n = 21   d_n = -0-1i 
assign X[4'b1110] [21] = 146'h 0000000000000000000000000000400000000;  // +0.0000000000000284 = 0.5 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+-1^2) * 2^(-2*22) )   n = 22   d_n = -0-1i 
assign X[4'b1110] [22] = 146'h 0000000000000000000000000000040000000;  // +0.0000000000000071 = 0.5 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+-1^2) * 2^(-2*23) )   n = 23   d_n = -0-1i 
assign X[4'b1110] [23] = 146'h 0000000000000000000000000000004000000;  // +0.0000000000000018 = 0.5 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+-1^2) * 2^(-2*24) )   n = 24   d_n = -0-1i 
assign X[4'b1110] [24] = 146'h 0000000000000000000000000000000400000;  // +0.0000000000000004 = 0.5 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+-1^2) * 2^(-2*25) )   n = 25   d_n = -0-1i 
assign X[4'b1110] [25] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+-1^2) * 2^(-2*26) )   n = 26   d_n = -0-1i 
assign X[4'b1110] [26] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+-1^2) * 2^(-2*27) )   n = 27   d_n = -0-1i 
assign X[4'b1110] [27] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+-1^2) * 2^(-2*28) )   n = 28   d_n = -0-1i 
assign X[4'b1110] [28] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+-1^2) * 2^(-2*29) )   n = 29   d_n = -0-1i 
assign X[4'b1110] [29] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+-1^2) * 2^(-2*30) )   n = 30   d_n = -0-1i 
assign X[4'b1110] [30] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+-1^2) * 2^(-2*31) )   n = 31   d_n = -0-1i 
assign X[4'b1110] [31] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+-1^2) * 2^(-2*32) )   n = 32   d_n = -0-1i 
assign X[4'b1110] [32] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+-1^2) * 2^(-2*33) )   n = 33   d_n = -0-1i 
assign X[4'b1110] [33] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+-1^2) * 2^(-2*34) )   n = 34   d_n = -0-1i 
assign X[4'b1110] [34] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+-1^2) * 2^(-2*35) )   n = 35   d_n = -0-1i 
assign X[4'b1110] [35] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+-1^2) * 2^(-2*36) )   n = 36   d_n = -0-1i 
assign X[4'b1110] [36] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+-1^2) * 2^(-2*37) )   n = 37   d_n = -0-1i 
assign X[4'b1110] [37] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+-1^2) * 2^(-2*38) )   n = 38   d_n = -0-1i 
assign X[4'b1110] [38] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+-1^2) * 2^(-2*39) )   n = 39   d_n = -0-1i 
assign X[4'b1110] [39] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+-1^2) * 2^(-2*40) )   n = 40   d_n = -0-1i 
assign X[4'b1110] [40] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+-1^2) * 2^(-2*41) )   n = 41   d_n = -0-1i 
assign X[4'b1110] [41] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+-1^2) * 2^(-2*42) )   n = 42   d_n = -0-1i 
assign X[4'b1110] [42] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+-1^2) * 2^(-2*43) )   n = 43   d_n = -0-1i 
assign X[4'b1110] [43] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+-1^2) * 2^(-2*44) )   n = 44   d_n = -0-1i 
assign X[4'b1110] [44] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+-1^2) * 2^(-2*45) )   n = 45   d_n = -0-1i 
assign X[4'b1110] [45] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+-1^2) * 2^(-2*46) )   n = 46   d_n = -0-1i 
assign X[4'b1110] [46] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+-1^2) * 2^(-2*47) )   n = 47   d_n = -0-1i 
assign X[4'b1110] [47] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+-1^2) * 2^(-2*48) )   n = 48   d_n = -0-1i 
assign X[4'b1110] [48] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+-1^2) * 2^(-2*49) )   n = 49   d_n = -0-1i 
assign X[4'b1110] [49] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+-1^2) * 2^(-2*50) )   n = 50   d_n = -0-1i 
assign X[4'b1110] [50] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+-1^2) * 2^(-2*51) )   n = 51   d_n = -0-1i 
assign X[4'b1110] [51] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+-1^2) * 2^(-2*52) )   n = 52   d_n = -0-1i 
assign X[4'b1110] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+-1^2) * 2^(-2*53) )   n = 53   d_n = -0-1i 
assign X[4'b1110] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+-1^2) * 2^(-2*54) )   n = 54   d_n = -0-1i 
assign X[4'b1110] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+-1^2) * 2^(-2*55) )   n = 55   d_n = -0-1i 
assign X[4'b1110] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+-1^2) * 2^(-2*56) )   n = 56   d_n = -0-1i 
assign X[4'b1110] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+-1^2) * 2^(-2*57) )   n = 57   d_n = -0-1i 
assign X[4'b1110] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+-1^2) * 2^(-2*58) )   n = 58   d_n = -0-1i 
assign X[4'b1110] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+-1^2) * 2^(-2*59) )   n = 59   d_n = -0-1i 
assign X[4'b1110] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+-1^2) * 2^(-2*60) )   n = 60   d_n = -0-1i 
assign X[4'b1110] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+-1^2) * 2^(-2*61) )   n = 61   d_n = -0-1i 
assign X[4'b1110] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+-1^2) * 2^(-2*62) )   n = 62   d_n = -0-1i 
assign X[4'b1110] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+-1^2) * 2^(-2*63) )   n = 63   d_n = -0-1i 
assign X[4'b1110] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+-1^2) * 2^(-2*64) )   n = 64   d_n = -0-1i 
assign X[4'b1111] [00] = 146'h 000000C443104303100000000000000000000;  // -0.3465735902799726 = 0.5 * ln( 1 + -1 * 2^(-1+1) + (-1^2+-1^2) * 2^(-2*1) )   n =  1   d_n = -1-1i 
assign X[4'b1111] [01] = 146'h 00000030100CC303303200000000000000000;  // -0.2350018146228677 = 0.5 * ln( 1 + -1 * 2^(-2+1) + (-1^2+-1^2) * 2^(-2*2) )   n =  2   d_n = -1-1i 
assign X[4'b1111] [02] = 146'h 0000000C004C430C10C100000000000000000;  // -0.1234300389657629 = 0.5 * ln( 1 + -1 * 2^(-3+1) + (-1^2+-1^2) * 2^(-2*3) )   n =  3   d_n = -1-1i 
assign X[4'b1111] [03] = 146'h 0000000300013030C0CC20000000000000000;  // -0.0623212226036383 = 0.5 * ln( 1 + -1 * 2^(-4+1) + (-1^2+-1^2) * 2^(-2*4) )   n =  4   d_n = -1-1i 
assign X[4'b1111] [04] = 146'h 00000000C00004CC4C3030000000000000000;  // -0.0312286774668733 = 0.5 * ln( 1 + -1 * 2^(-5+1) + (-1^2+-1^2) * 2^(-2*5) )   n =  5   d_n = -1-1i 
assign X[4'b1111] [05] = 146'h 000000003000001330330C000000000000000;  // -0.0156223965190538 = 0.5 * ln( 1 + -1 * 2^(-6+1) + (-1^2+-1^2) * 2^(-2*6) )   n =  6   d_n = -1-1i 
assign X[4'b1111] [06] = 146'h 000000000C0000004CCC4D000000000000000;  // -0.0078121783599899 = 0.5 * ln( 1 + -1 * 2^(-7+1) + (-1^2+-1^2) * 2^(-2*7) )   n =  7   d_n = -1-1i 
assign X[4'b1111] [07] = 146'h 0000000003000000013330400000000000000;  // -0.0039062100300119 = 0.5 * ln( 1 + -1 * 2^(-8+1) + (-1^2+-1^2) * 2^(-2*8) )   n =  8   d_n = -1-1i 
assign X[4'b1111] [08] = 146'h 0000000000C000000004CCD00000000000000;  // -0.0019531200183716 = 0.5 * ln( 1 + -1 * 2^(-9+1) + (-1^2+-1^2) * 2^(-2*9) )   n =  9   d_n = -1-1i 
assign X[4'b1111] [09] = 146'h 0000000000300000000013340000000000000;  // -0.0009765618782081 = 0.5 * ln( 1 + -1 * 2^(-10+1) + (-1^2+-1^2) * 2^(-2*10) )   n = 10   d_n = -1-1i 
assign X[4'b1111] [10] = 146'h 00000000000C00000000004D0000000000000;  // -0.0004882811723329 = 0.5 * ln( 1 + -1 * 2^(-11+1) + (-1^2+-1^2) * 2^(-2*11) )   n = 11   d_n = -1-1i 
assign X[4'b1111] [11] = 146'h 0000000000030000000000014000000000000;  // -0.0002441406152952 = 0.5 * ln( 1 + -1 * 2^(-12+1) + (-1^2+-1^2) * 2^(-2*12) )   n = 12   d_n = -1-1i 
assign X[4'b1111] [12] = 146'h 000000000000C000000000000800000000000;  // -0.0001220703112871 = 0.5 * ln( 1 + -1 * 2^(-13+1) + (-1^2+-1^2) * 2^(-2*13) )   n = 13   d_n = -1-1i 
assign X[4'b1111] [13] = 146'h 0000000000003000000000000000000000000;  // -0.0000610351560984 = 0.5 * ln( 1 + -1 * 2^(-14+1) + (-1^2+-1^2) * 2^(-2*14) )   n = 14   d_n = -1-1i 
assign X[4'b1111] [14] = 146'h 0000000000000C00000000000000000000000;  // -0.0000305175781061 = 0.5 * ln( 1 + -1 * 2^(-15+1) + (-1^2+-1^2) * 2^(-2*15) )   n = 15   d_n = -1-1i 
assign X[4'b1111] [15] = 146'h 0000000000000300000000000000000000000;  // -0.0000152587890601 = 0.5 * ln( 1 + -1 * 2^(-16+1) + (-1^2+-1^2) * 2^(-2*16) )   n = 16   d_n = -1-1i 
assign X[4'b1111] [16] = 146'h 00000000000000C0000000000000000000000;  // -0.0000076293945310 = 0.5 * ln( 1 + -1 * 2^(-17+1) + (-1^2+-1^2) * 2^(-2*17) )   n = 17   d_n = -1-1i 
assign X[4'b1111] [17] = 146'h 0000000000000030000000000000000000000;  // -0.0000038146972656 = 0.5 * ln( 1 + -1 * 2^(-18+1) + (-1^2+-1^2) * 2^(-2*18) )   n = 18   d_n = -1-1i 
assign X[4'b1111] [18] = 146'h 000000000000000C000000000000000000000;  // -0.0000019073486328 = 0.5 * ln( 1 + -1 * 2^(-19+1) + (-1^2+-1^2) * 2^(-2*19) )   n = 19   d_n = -1-1i 
assign X[4'b1111] [19] = 146'h 0000000000000003000000000000000000000;  // -0.0000009536743164 = 0.5 * ln( 1 + -1 * 2^(-20+1) + (-1^2+-1^2) * 2^(-2*20) )   n = 20   d_n = -1-1i 
assign X[4'b1111] [20] = 146'h 0000000000000000C00000000000000000000;  // -0.0000004768371582 = 0.5 * ln( 1 + -1 * 2^(-21+1) + (-1^2+-1^2) * 2^(-2*21) )   n = 21   d_n = -1-1i 
assign X[4'b1111] [21] = 146'h 0000000000000000300000000000000000000;  // -0.0000002384185791 = 0.5 * ln( 1 + -1 * 2^(-22+1) + (-1^2+-1^2) * 2^(-2*22) )   n = 22   d_n = -1-1i 
assign X[4'b1111] [22] = 146'h 00000000000000000C0000000000000000000;  // -0.0000001192092896 = 0.5 * ln( 1 + -1 * 2^(-23+1) + (-1^2+-1^2) * 2^(-2*23) )   n = 23   d_n = -1-1i 
assign X[4'b1111] [23] = 146'h 0000000000000000030000000000000000000;  // -0.0000000596046448 = 0.5 * ln( 1 + -1 * 2^(-24+1) + (-1^2+-1^2) * 2^(-2*24) )   n = 24   d_n = -1-1i 
assign X[4'b1111] [24] = 146'h 000000000000000000C000000000000000000;  // -0.0000000298023224 = 0.5 * ln( 1 + -1 * 2^(-25+1) + (-1^2+-1^2) * 2^(-2*25) )   n = 25   d_n = -1-1i 
assign X[4'b1111] [25] = 146'h 0000000000000000003000000000000000000;  // -0.0000000149011612 = 0.5 * ln( 1 + -1 * 2^(-26+1) + (-1^2+-1^2) * 2^(-2*26) )   n = 26   d_n = -1-1i 
assign X[4'b1111] [26] = 146'h 0000000000000000000C00000000000000000;  // -0.0000000074505806 = 0.5 * ln( 1 + -1 * 2^(-27+1) + (-1^2+-1^2) * 2^(-2*27) )   n = 27   d_n = -1-1i 
assign X[4'b1111] [27] = 146'h 0000000000000000000300000000000000000;  // -0.0000000037252903 = 0.5 * ln( 1 + -1 * 2^(-28+1) + (-1^2+-1^2) * 2^(-2*28) )   n = 28   d_n = -1-1i 
assign X[4'b1111] [28] = 146'h 00000000000000000000C0000000000000000;  // -0.0000000018626452 = 0.5 * ln( 1 + -1 * 2^(-29+1) + (-1^2+-1^2) * 2^(-2*29) )   n = 29   d_n = -1-1i 
assign X[4'b1111] [29] = 146'h 0000000000000000000030000000000000000;  // -0.0000000009313226 = 0.5 * ln( 1 + -1 * 2^(-30+1) + (-1^2+-1^2) * 2^(-2*30) )   n = 30   d_n = -1-1i 
assign X[4'b1111] [30] = 146'h 000000000000000000000C000000000000000;  // -0.0000000004656613 = 0.5 * ln( 1 + -1 * 2^(-31+1) + (-1^2+-1^2) * 2^(-2*31) )   n = 31   d_n = -1-1i 
assign X[4'b1111] [31] = 146'h 0000000000000000000003000000000000000;  // -0.0000000002328306 = 0.5 * ln( 1 + -1 * 2^(-32+1) + (-1^2+-1^2) * 2^(-2*32) )   n = 32   d_n = -1-1i 
assign X[4'b1111] [32] = 146'h 0000000000000000000000C00000000000000;  // -0.0000000001164153 = 0.5 * ln( 1 + -1 * 2^(-33+1) + (-1^2+-1^2) * 2^(-2*33) )   n = 33   d_n = -1-1i 
assign X[4'b1111] [33] = 146'h 0000000000000000000000300000000000000;  // -0.0000000000582077 = 0.5 * ln( 1 + -1 * 2^(-34+1) + (-1^2+-1^2) * 2^(-2*34) )   n = 34   d_n = -1-1i 
assign X[4'b1111] [34] = 146'h 00000000000000000000000C0000000000000;  // -0.0000000000291038 = 0.5 * ln( 1 + -1 * 2^(-35+1) + (-1^2+-1^2) * 2^(-2*35) )   n = 35   d_n = -1-1i 
assign X[4'b1111] [35] = 146'h 0000000000000000000000030000000000000;  // -0.0000000000145519 = 0.5 * ln( 1 + -1 * 2^(-36+1) + (-1^2+-1^2) * 2^(-2*36) )   n = 36   d_n = -1-1i 
assign X[4'b1111] [36] = 146'h 000000000000000000000000C000000000000;  // -0.0000000000072760 = 0.5 * ln( 1 + -1 * 2^(-37+1) + (-1^2+-1^2) * 2^(-2*37) )   n = 37   d_n = -1-1i 
assign X[4'b1111] [37] = 146'h 0000000000000000000000003000000000000;  // -0.0000000000036380 = 0.5 * ln( 1 + -1 * 2^(-38+1) + (-1^2+-1^2) * 2^(-2*38) )   n = 38   d_n = -1-1i 
assign X[4'b1111] [38] = 146'h 0000000000000000000000000C00000000000;  // -0.0000000000018190 = 0.5 * ln( 1 + -1 * 2^(-39+1) + (-1^2+-1^2) * 2^(-2*39) )   n = 39   d_n = -1-1i 
assign X[4'b1111] [39] = 146'h 0000000000000000000000000300000000000;  // -0.0000000000009095 = 0.5 * ln( 1 + -1 * 2^(-40+1) + (-1^2+-1^2) * 2^(-2*40) )   n = 40   d_n = -1-1i 
assign X[4'b1111] [40] = 146'h 00000000000000000000000000C0000000000;  // -0.0000000000004547 = 0.5 * ln( 1 + -1 * 2^(-41+1) + (-1^2+-1^2) * 2^(-2*41) )   n = 41   d_n = -1-1i 
assign X[4'b1111] [41] = 146'h 0000000000000000000000000030000000000;  // -0.0000000000002274 = 0.5 * ln( 1 + -1 * 2^(-42+1) + (-1^2+-1^2) * 2^(-2*42) )   n = 42   d_n = -1-1i 
assign X[4'b1111] [42] = 146'h 000000000000000000000000000C000000000;  // -0.0000000000001137 = 0.5 * ln( 1 + -1 * 2^(-43+1) + (-1^2+-1^2) * 2^(-2*43) )   n = 43   d_n = -1-1i 
assign X[4'b1111] [43] = 146'h 0000000000000000000000000003000000000;  // -0.0000000000000568 = 0.5 * ln( 1 + -1 * 2^(-44+1) + (-1^2+-1^2) * 2^(-2*44) )   n = 44   d_n = -1-1i 
assign X[4'b1111] [44] = 146'h 0000000000000000000000000000C00000000;  // -0.0000000000000284 = 0.5 * ln( 1 + -1 * 2^(-45+1) + (-1^2+-1^2) * 2^(-2*45) )   n = 45   d_n = -1-1i 
assign X[4'b1111] [45] = 146'h 0000000000000000000000000000300000000;  // -0.0000000000000142 = 0.5 * ln( 1 + -1 * 2^(-46+1) + (-1^2+-1^2) * 2^(-2*46) )   n = 46   d_n = -1-1i 
assign X[4'b1111] [46] = 146'h 00000000000000000000000000000C0000000;  // -0.0000000000000071 = 0.5 * ln( 1 + -1 * 2^(-47+1) + (-1^2+-1^2) * 2^(-2*47) )   n = 47   d_n = -1-1i 
assign X[4'b1111] [47] = 146'h 0000000000000000000000000000030000000;  // -0.0000000000000036 = 0.5 * ln( 1 + -1 * 2^(-48+1) + (-1^2+-1^2) * 2^(-2*48) )   n = 48   d_n = -1-1i 
assign X[4'b1111] [48] = 146'h 000000000000000000000000000000C000000;  // -0.0000000000000018 = 0.5 * ln( 1 + -1 * 2^(-49+1) + (-1^2+-1^2) * 2^(-2*49) )   n = 49   d_n = -1-1i 
assign X[4'b1111] [49] = 146'h 0000000000000000000000000000003000000;  // -0.0000000000000009 = 0.5 * ln( 1 + -1 * 2^(-50+1) + (-1^2+-1^2) * 2^(-2*50) )   n = 50   d_n = -1-1i 
assign X[4'b1111] [50] = 146'h 0000000000000000000000000000000C00000;  // -0.0000000000000004 = 0.5 * ln( 1 + -1 * 2^(-51+1) + (-1^2+-1^2) * 2^(-2*51) )   n = 51   d_n = -1-1i 
assign X[4'b1111] [51] = 146'h 0000000000000000000000000000000300000;  // -0.0000000000000002 = 0.5 * ln( 1 + -1 * 2^(-52+1) + (-1^2+-1^2) * 2^(-2*52) )   n = 52   d_n = -1-1i 
assign X[4'b1111] [52] = 146'h 00000000000000000000000000000000C0000;  // -0.0000000000000001 = 0.5 * ln( 1 + -1 * 2^(-53+1) + (-1^2+-1^2) * 2^(-2*53) )   n = 53   d_n = -1-1i 
assign X[4'b1111] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-54+1) + (-1^2+-1^2) * 2^(-2*54) )   n = 54   d_n = -1-1i 
assign X[4'b1111] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-55+1) + (-1^2+-1^2) * 2^(-2*55) )   n = 55   d_n = -1-1i 
assign X[4'b1111] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-56+1) + (-1^2+-1^2) * 2^(-2*56) )   n = 56   d_n = -1-1i 
assign X[4'b1111] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-57+1) + (-1^2+-1^2) * 2^(-2*57) )   n = 57   d_n = -1-1i 
assign X[4'b1111] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-58+1) + (-1^2+-1^2) * 2^(-2*58) )   n = 58   d_n = -1-1i 
assign X[4'b1111] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-59+1) + (-1^2+-1^2) * 2^(-2*59) )   n = 59   d_n = -1-1i 
assign X[4'b1111] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-60+1) + (-1^2+-1^2) * 2^(-2*60) )   n = 60   d_n = -1-1i 
assign X[4'b1111] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-61+1) + (-1^2+-1^2) * 2^(-2*61) )   n = 61   d_n = -1-1i 
assign X[4'b1111] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-62+1) + (-1^2+-1^2) * 2^(-2*62) )   n = 62   d_n = -1-1i 
assign X[4'b1111] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-63+1) + (-1^2+-1^2) * 2^(-2*63) )   n = 63   d_n = -1-1i 
assign X[4'b1111] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-64+1) + (-1^2+-1^2) * 2^(-2*64) )   n = 64   d_n = -1-1i 
assign Y[4'b0000] [00] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = 0 
assign Y[4'b0000] [01] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = 0 
assign Y[4'b0000] [02] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = 0 
assign Y[4'b0000] [03] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = 0 
assign Y[4'b0000] [04] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = 0 
assign Y[4'b0000] [05] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = 0 
assign Y[4'b0000] [06] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = 0 
assign Y[4'b0000] [07] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = 0 
assign Y[4'b0000] [08] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = 0 
assign Y[4'b0000] [09] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = 0 
assign Y[4'b0000] [10] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = 0 
assign Y[4'b0000] [11] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = 0 
assign Y[4'b0000] [12] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = 0 
assign Y[4'b0000] [13] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = 0 
assign Y[4'b0000] [14] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = 0 
assign Y[4'b0000] [15] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = 0 
assign Y[4'b0000] [16] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = 0 
assign Y[4'b0000] [17] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = 0 
assign Y[4'b0000] [18] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = 0 
assign Y[4'b0000] [19] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = 0 
assign Y[4'b0000] [20] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = 0 
assign Y[4'b0000] [21] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = 0 
assign Y[4'b0000] [22] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = 0 
assign Y[4'b0000] [23] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = 0 
assign Y[4'b0000] [24] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = 0 
assign Y[4'b0000] [25] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = 0 
assign Y[4'b0000] [26] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = 0 
assign Y[4'b0000] [27] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = 0 
assign Y[4'b0000] [28] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = 0 
assign Y[4'b0000] [29] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = 0 
assign Y[4'b0000] [30] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = 0 
assign Y[4'b0000] [31] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = 0 
assign Y[4'b0000] [32] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = 0 
assign Y[4'b0000] [33] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = 0 
assign Y[4'b0000] [34] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = 0 
assign Y[4'b0000] [35] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = 0 
assign Y[4'b0000] [36] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = 0 
assign Y[4'b0000] [37] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = 0 
assign Y[4'b0000] [38] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = 0 
assign Y[4'b0000] [39] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = 0 
assign Y[4'b0000] [40] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = 0 
assign Y[4'b0000] [41] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = 0 
assign Y[4'b0000] [42] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = 0 
assign Y[4'b0000] [43] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = 0 
assign Y[4'b0000] [44] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = 0 
assign Y[4'b0000] [45] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = 0 
assign Y[4'b0000] [46] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = 0 
assign Y[4'b0000] [47] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = 0 
assign Y[4'b0000] [48] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = 0 
assign Y[4'b0000] [49] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = 0 
assign Y[4'b0000] [50] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = 0 
assign Y[4'b0000] [51] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = 0 
assign Y[4'b0000] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = 0 
assign Y[4'b0000] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = 0 
assign Y[4'b0000] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = 0 
assign Y[4'b0000] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = 0 
assign Y[4'b0000] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = 0 
assign Y[4'b0000] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = 0 
assign Y[4'b0000] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = 0 
assign Y[4'b0000] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = 0 
assign Y[4'b0000] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = 0 
assign Y[4'b0000] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = 0 
assign Y[4'b0000] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = 0 
assign Y[4'b0000] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = 0 
assign Y[4'b0001] [00] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^1 ) )   n =  1   d_n = 1 
assign Y[4'b0001] [01] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^2 ) )   n =  2   d_n = 1 
assign Y[4'b0001] [02] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^3 ) )   n =  3   d_n = 1 
assign Y[4'b0001] [03] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^4 ) )   n =  4   d_n = 1 
assign Y[4'b0001] [04] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^5 ) )   n =  5   d_n = 1 
assign Y[4'b0001] [05] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^6 ) )   n =  6   d_n = 1 
assign Y[4'b0001] [06] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^7 ) )   n =  7   d_n = 1 
assign Y[4'b0001] [07] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^8 ) )   n =  8   d_n = 1 
assign Y[4'b0001] [08] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^9 ) )   n =  9   d_n = 1 
assign Y[4'b0001] [09] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^10 ) )   n = 10   d_n = 1 
assign Y[4'b0001] [10] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^11 ) )   n = 11   d_n = 1 
assign Y[4'b0001] [11] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^12 ) )   n = 12   d_n = 1 
assign Y[4'b0001] [12] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^13 ) )   n = 13   d_n = 1 
assign Y[4'b0001] [13] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^14 ) )   n = 14   d_n = 1 
assign Y[4'b0001] [14] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^15 ) )   n = 15   d_n = 1 
assign Y[4'b0001] [15] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^16 ) )   n = 16   d_n = 1 
assign Y[4'b0001] [16] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^17 ) )   n = 17   d_n = 1 
assign Y[4'b0001] [17] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^18 ) )   n = 18   d_n = 1 
assign Y[4'b0001] [18] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^19 ) )   n = 19   d_n = 1 
assign Y[4'b0001] [19] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^20 ) )   n = 20   d_n = 1 
assign Y[4'b0001] [20] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^21 ) )   n = 21   d_n = 1 
assign Y[4'b0001] [21] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^22 ) )   n = 22   d_n = 1 
assign Y[4'b0001] [22] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^23 ) )   n = 23   d_n = 1 
assign Y[4'b0001] [23] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^24 ) )   n = 24   d_n = 1 
assign Y[4'b0001] [24] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^25 ) )   n = 25   d_n = 1 
assign Y[4'b0001] [25] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^26 ) )   n = 26   d_n = 1 
assign Y[4'b0001] [26] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^27 ) )   n = 27   d_n = 1 
assign Y[4'b0001] [27] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^28 ) )   n = 28   d_n = 1 
assign Y[4'b0001] [28] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^29 ) )   n = 29   d_n = 1 
assign Y[4'b0001] [29] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^30 ) )   n = 30   d_n = 1 
assign Y[4'b0001] [30] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^31 ) )   n = 31   d_n = 1 
assign Y[4'b0001] [31] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^32 ) )   n = 32   d_n = 1 
assign Y[4'b0001] [32] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^33 ) )   n = 33   d_n = 1 
assign Y[4'b0001] [33] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^34 ) )   n = 34   d_n = 1 
assign Y[4'b0001] [34] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^35 ) )   n = 35   d_n = 1 
assign Y[4'b0001] [35] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^36 ) )   n = 36   d_n = 1 
assign Y[4'b0001] [36] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^37 ) )   n = 37   d_n = 1 
assign Y[4'b0001] [37] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^38 ) )   n = 38   d_n = 1 
assign Y[4'b0001] [38] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^39 ) )   n = 39   d_n = 1 
assign Y[4'b0001] [39] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^40 ) )   n = 40   d_n = 1 
assign Y[4'b0001] [40] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^41 ) )   n = 41   d_n = 1 
assign Y[4'b0001] [41] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^42 ) )   n = 42   d_n = 1 
assign Y[4'b0001] [42] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^43 ) )   n = 43   d_n = 1 
assign Y[4'b0001] [43] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^44 ) )   n = 44   d_n = 1 
assign Y[4'b0001] [44] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^45 ) )   n = 45   d_n = 1 
assign Y[4'b0001] [45] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^46 ) )   n = 46   d_n = 1 
assign Y[4'b0001] [46] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^47 ) )   n = 47   d_n = 1 
assign Y[4'b0001] [47] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^48 ) )   n = 48   d_n = 1 
assign Y[4'b0001] [48] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^49 ) )   n = 49   d_n = 1 
assign Y[4'b0001] [49] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^50 ) )   n = 50   d_n = 1 
assign Y[4'b0001] [50] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^51 ) )   n = 51   d_n = 1 
assign Y[4'b0001] [51] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^52 ) )   n = 52   d_n = 1 
assign Y[4'b0001] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^53 ) )   n = 53   d_n = 1 
assign Y[4'b0001] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^54 ) )   n = 54   d_n = 1 
assign Y[4'b0001] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^55 ) )   n = 55   d_n = 1 
assign Y[4'b0001] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^56 ) )   n = 56   d_n = 1 
assign Y[4'b0001] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^57 ) )   n = 57   d_n = 1 
assign Y[4'b0001] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^58 ) )   n = 58   d_n = 1 
assign Y[4'b0001] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^59 ) )   n = 59   d_n = 1 
assign Y[4'b0001] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^60 ) )   n = 60   d_n = 1 
assign Y[4'b0001] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^61 ) )   n = 61   d_n = 1 
assign Y[4'b0001] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^62 ) )   n = 62   d_n = 1 
assign Y[4'b0001] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^63 ) )   n = 63   d_n = 1 
assign Y[4'b0001] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^64 ) )   n = 64   d_n = 1 
assign Y[4'b0010] [00] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = -0 
assign Y[4'b0010] [01] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = -0 
assign Y[4'b0010] [02] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = -0 
assign Y[4'b0010] [03] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = -0 
assign Y[4'b0010] [04] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = -0 
assign Y[4'b0010] [05] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = -0 
assign Y[4'b0010] [06] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = -0 
assign Y[4'b0010] [07] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = -0 
assign Y[4'b0010] [08] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = -0 
assign Y[4'b0010] [09] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = -0 
assign Y[4'b0010] [10] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = -0 
assign Y[4'b0010] [11] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = -0 
assign Y[4'b0010] [12] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = -0 
assign Y[4'b0010] [13] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = -0 
assign Y[4'b0010] [14] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = -0 
assign Y[4'b0010] [15] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = -0 
assign Y[4'b0010] [16] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = -0 
assign Y[4'b0010] [17] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = -0 
assign Y[4'b0010] [18] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = -0 
assign Y[4'b0010] [19] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = -0 
assign Y[4'b0010] [20] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = -0 
assign Y[4'b0010] [21] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = -0 
assign Y[4'b0010] [22] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = -0 
assign Y[4'b0010] [23] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = -0 
assign Y[4'b0010] [24] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = -0 
assign Y[4'b0010] [25] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = -0 
assign Y[4'b0010] [26] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = -0 
assign Y[4'b0010] [27] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = -0 
assign Y[4'b0010] [28] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = -0 
assign Y[4'b0010] [29] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = -0 
assign Y[4'b0010] [30] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = -0 
assign Y[4'b0010] [31] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = -0 
assign Y[4'b0010] [32] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = -0 
assign Y[4'b0010] [33] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = -0 
assign Y[4'b0010] [34] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = -0 
assign Y[4'b0010] [35] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = -0 
assign Y[4'b0010] [36] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = -0 
assign Y[4'b0010] [37] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = -0 
assign Y[4'b0010] [38] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = -0 
assign Y[4'b0010] [39] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = -0 
assign Y[4'b0010] [40] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = -0 
assign Y[4'b0010] [41] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = -0 
assign Y[4'b0010] [42] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = -0 
assign Y[4'b0010] [43] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = -0 
assign Y[4'b0010] [44] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = -0 
assign Y[4'b0010] [45] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = -0 
assign Y[4'b0010] [46] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = -0 
assign Y[4'b0010] [47] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = -0 
assign Y[4'b0010] [48] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = -0 
assign Y[4'b0010] [49] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = -0 
assign Y[4'b0010] [50] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = -0 
assign Y[4'b0010] [51] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = -0 
assign Y[4'b0010] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = -0 
assign Y[4'b0010] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = -0 
assign Y[4'b0010] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = -0 
assign Y[4'b0010] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = -0 
assign Y[4'b0010] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = -0 
assign Y[4'b0010] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = -0 
assign Y[4'b0010] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = -0 
assign Y[4'b0010] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = -0 
assign Y[4'b0010] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = -0 
assign Y[4'b0010] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = -0 
assign Y[4'b0010] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = -0 
assign Y[4'b0010] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = -0 
assign Y[4'b0011] [00] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^1 ) )   n =  1   d_n = -1 
assign Y[4'b0011] [01] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^2 ) )   n =  2   d_n = -1 
assign Y[4'b0011] [02] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^3 ) )   n =  3   d_n = -1 
assign Y[4'b0011] [03] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^4 ) )   n =  4   d_n = -1 
assign Y[4'b0011] [04] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^5 ) )   n =  5   d_n = -1 
assign Y[4'b0011] [05] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^6 ) )   n =  6   d_n = -1 
assign Y[4'b0011] [06] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^7 ) )   n =  7   d_n = -1 
assign Y[4'b0011] [07] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^8 ) )   n =  8   d_n = -1 
assign Y[4'b0011] [08] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^9 ) )   n =  9   d_n = -1 
assign Y[4'b0011] [09] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^10 ) )   n = 10   d_n = -1 
assign Y[4'b0011] [10] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^11 ) )   n = 11   d_n = -1 
assign Y[4'b0011] [11] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^12 ) )   n = 12   d_n = -1 
assign Y[4'b0011] [12] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^13 ) )   n = 13   d_n = -1 
assign Y[4'b0011] [13] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^14 ) )   n = 14   d_n = -1 
assign Y[4'b0011] [14] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^15 ) )   n = 15   d_n = -1 
assign Y[4'b0011] [15] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^16 ) )   n = 16   d_n = -1 
assign Y[4'b0011] [16] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^17 ) )   n = 17   d_n = -1 
assign Y[4'b0011] [17] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^18 ) )   n = 18   d_n = -1 
assign Y[4'b0011] [18] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^19 ) )   n = 19   d_n = -1 
assign Y[4'b0011] [19] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^20 ) )   n = 20   d_n = -1 
assign Y[4'b0011] [20] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^21 ) )   n = 21   d_n = -1 
assign Y[4'b0011] [21] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^22 ) )   n = 22   d_n = -1 
assign Y[4'b0011] [22] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^23 ) )   n = 23   d_n = -1 
assign Y[4'b0011] [23] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^24 ) )   n = 24   d_n = -1 
assign Y[4'b0011] [24] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^25 ) )   n = 25   d_n = -1 
assign Y[4'b0011] [25] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^26 ) )   n = 26   d_n = -1 
assign Y[4'b0011] [26] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^27 ) )   n = 27   d_n = -1 
assign Y[4'b0011] [27] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^28 ) )   n = 28   d_n = -1 
assign Y[4'b0011] [28] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^29 ) )   n = 29   d_n = -1 
assign Y[4'b0011] [29] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^30 ) )   n = 30   d_n = -1 
assign Y[4'b0011] [30] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^31 ) )   n = 31   d_n = -1 
assign Y[4'b0011] [31] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^32 ) )   n = 32   d_n = -1 
assign Y[4'b0011] [32] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^33 ) )   n = 33   d_n = -1 
assign Y[4'b0011] [33] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^34 ) )   n = 34   d_n = -1 
assign Y[4'b0011] [34] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^35 ) )   n = 35   d_n = -1 
assign Y[4'b0011] [35] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^36 ) )   n = 36   d_n = -1 
assign Y[4'b0011] [36] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^37 ) )   n = 37   d_n = -1 
assign Y[4'b0011] [37] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^38 ) )   n = 38   d_n = -1 
assign Y[4'b0011] [38] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^39 ) )   n = 39   d_n = -1 
assign Y[4'b0011] [39] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^40 ) )   n = 40   d_n = -1 
assign Y[4'b0011] [40] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^41 ) )   n = 41   d_n = -1 
assign Y[4'b0011] [41] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^42 ) )   n = 42   d_n = -1 
assign Y[4'b0011] [42] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^43 ) )   n = 43   d_n = -1 
assign Y[4'b0011] [43] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^44 ) )   n = 44   d_n = -1 
assign Y[4'b0011] [44] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^45 ) )   n = 45   d_n = -1 
assign Y[4'b0011] [45] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^46 ) )   n = 46   d_n = -1 
assign Y[4'b0011] [46] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^47 ) )   n = 47   d_n = -1 
assign Y[4'b0011] [47] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^48 ) )   n = 48   d_n = -1 
assign Y[4'b0011] [48] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^49 ) )   n = 49   d_n = -1 
assign Y[4'b0011] [49] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^50 ) )   n = 50   d_n = -1 
assign Y[4'b0011] [50] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^51 ) )   n = 51   d_n = -1 
assign Y[4'b0011] [51] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^52 ) )   n = 52   d_n = -1 
assign Y[4'b0011] [52] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^53 ) )   n = 53   d_n = -1 
assign Y[4'b0011] [53] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^54 ) )   n = 54   d_n = -1 
assign Y[4'b0011] [54] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^55 ) )   n = 55   d_n = -1 
assign Y[4'b0011] [55] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^56 ) )   n = 56   d_n = -1 
assign Y[4'b0011] [56] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^57 ) )   n = 57   d_n = -1 
assign Y[4'b0011] [57] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^58 ) )   n = 58   d_n = -1 
assign Y[4'b0011] [58] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^59 ) )   n = 59   d_n = -1 
assign Y[4'b0011] [59] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^60 ) )   n = 60   d_n = -1 
assign Y[4'b0011] [60] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^61 ) )   n = 61   d_n = -1 
assign Y[4'b0011] [61] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^62 ) )   n = 62   d_n = -1 
assign Y[4'b0011] [62] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^63 ) )   n = 63   d_n = -1 
assign Y[4'b0011] [63] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^64 ) )   n = 64   d_n = -1 
assign Y[4'b0100] [00] = 146'h 00000040C33304C4300400000000000000000;  // +0.4636476090008061 =  1 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = 0+1i 
assign Y[4'b0100] [01] = 146'h 000000100330C303300300000000000000000;  // +0.2449786631268641 =  1 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = 0+1i 
assign Y[4'b0100] [02] = 146'h 00000004000CCC30C44440000000000000000;  // +0.1243549945467614 =  1 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = 0+1i 
assign Y[4'b0100] [03] = 146'h 00000001000033330C0C30000000000000000;  // +0.0624188099959574 =  1 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = 0+1i 
assign Y[4'b0100] [04] = 146'h 00000000400000CCCCC304000000000000000;  // +0.0312398334302683 =  1 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = 0+1i 
assign Y[4'b0100] [05] = 146'h 0000000010000003333331000000000000000;  // +0.0156237286204768 =  1 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = 0+1i 
assign Y[4'b0100] [06] = 146'h 00000000040000000CCCCCC00000000000000;  // +0.0078123410601011 =  1 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = 0+1i 
assign Y[4'b0100] [07] = 146'h 0000000001000000003333300000000000000;  // +0.0039062301319670 =  1 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = 0+1i 
assign Y[4'b0100] [08] = 146'h 00000000004000000000CCCC0000000000000;  // +0.0019531225164788 =  1 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = 0+1i 
assign Y[4'b0100] [09] = 146'h 0000000000100000000003330000000000000;  // +0.0009765621895593 =  1 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = 0+1i 
assign Y[4'b0100] [10] = 146'h 00000000000400000000000CC000000000000;  // +0.0004882812111949 =  1 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = 0+1i 
assign Y[4'b0100] [11] = 146'h 0000000000010000000000003000000000000;  // +0.0002441406201494 =  1 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = 0+1i 
assign Y[4'b0100] [12] = 146'h 0000000000004000000000000400000000000;  // +0.0001220703118937 =  1 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = 0+1i 
assign Y[4'b0100] [13] = 146'h 0000000000001000000000000000000000000;  // +0.0000610351561742 =  1 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = 0+1i 
assign Y[4'b0100] [14] = 146'h 0000000000000400000000000000000000000;  // +0.0000305175781155 =  1 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = 0+1i 
assign Y[4'b0100] [15] = 146'h 0000000000000100000000000000000000000;  // +0.0000152587890613 =  1 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = 0+1i 
assign Y[4'b0100] [16] = 146'h 0000000000000040000000000000000000000;  // +0.0000076293945311 =  1 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = 0+1i 
assign Y[4'b0100] [17] = 146'h 0000000000000010000000000000000000000;  // +0.0000038146972656 =  1 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = 0+1i 
assign Y[4'b0100] [18] = 146'h 0000000000000004000000000000000000000;  // +0.0000019073486328 =  1 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = 0+1i 
assign Y[4'b0100] [19] = 146'h 0000000000000001000000000000000000000;  // +0.0000009536743164 =  1 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = 0+1i 
assign Y[4'b0100] [20] = 146'h 0000000000000000400000000000000000000;  // +0.0000004768371582 =  1 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = 0+1i 
assign Y[4'b0100] [21] = 146'h 0000000000000000100000000000000000000;  // +0.0000002384185791 =  1 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = 0+1i 
assign Y[4'b0100] [22] = 146'h 0000000000000000040000000000000000000;  // +0.0000001192092896 =  1 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = 0+1i 
assign Y[4'b0100] [23] = 146'h 0000000000000000010000000000000000000;  // +0.0000000596046448 =  1 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = 0+1i 
assign Y[4'b0100] [24] = 146'h 0000000000000000004000000000000000000;  // +0.0000000298023224 =  1 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = 0+1i 
assign Y[4'b0100] [25] = 146'h 0000000000000000001000000000000000000;  // +0.0000000149011612 =  1 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = 0+1i 
assign Y[4'b0100] [26] = 146'h 0000000000000000000400000000000000000;  // +0.0000000074505806 =  1 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = 0+1i 
assign Y[4'b0100] [27] = 146'h 0000000000000000000100000000000000000;  // +0.0000000037252903 =  1 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = 0+1i 
assign Y[4'b0100] [28] = 146'h 0000000000000000000040000000000000000;  // +0.0000000018626451 =  1 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = 0+1i 
assign Y[4'b0100] [29] = 146'h 0000000000000000000010000000000000000;  // +0.0000000009313226 =  1 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = 0+1i 
assign Y[4'b0100] [30] = 146'h 0000000000000000000004000000000000000;  // +0.0000000004656613 =  1 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = 0+1i 
assign Y[4'b0100] [31] = 146'h 0000000000000000000001000000000000000;  // +0.0000000002328306 =  1 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = 0+1i 
assign Y[4'b0100] [32] = 146'h 0000000000000000000000400000000000000;  // +0.0000000001164153 =  1 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = 0+1i 
assign Y[4'b0100] [33] = 146'h 0000000000000000000000100000000000000;  // +0.0000000000582077 =  1 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = 0+1i 
assign Y[4'b0100] [34] = 146'h 0000000000000000000000040000000000000;  // +0.0000000000291038 =  1 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = 0+1i 
assign Y[4'b0100] [35] = 146'h 0000000000000000000000010000000000000;  // +0.0000000000145519 =  1 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = 0+1i 
assign Y[4'b0100] [36] = 146'h 0000000000000000000000004000000000000;  // +0.0000000000072760 =  1 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = 0+1i 
assign Y[4'b0100] [37] = 146'h 0000000000000000000000001000000000000;  // +0.0000000000036380 =  1 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = 0+1i 
assign Y[4'b0100] [38] = 146'h 0000000000000000000000000400000000000;  // +0.0000000000018190 =  1 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = 0+1i 
assign Y[4'b0100] [39] = 146'h 0000000000000000000000000100000000000;  // +0.0000000000009095 =  1 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = 0+1i 
assign Y[4'b0100] [40] = 146'h 0000000000000000000000000040000000000;  // +0.0000000000004547 =  1 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = 0+1i 
assign Y[4'b0100] [41] = 146'h 0000000000000000000000000010000000000;  // +0.0000000000002274 =  1 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = 0+1i 
assign Y[4'b0100] [42] = 146'h 0000000000000000000000000004000000000;  // +0.0000000000001137 =  1 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = 0+1i 
assign Y[4'b0100] [43] = 146'h 0000000000000000000000000001000000000;  // +0.0000000000000568 =  1 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = 0+1i 
assign Y[4'b0100] [44] = 146'h 0000000000000000000000000000400000000;  // +0.0000000000000284 =  1 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = 0+1i 
assign Y[4'b0100] [45] = 146'h 0000000000000000000000000000100000000;  // +0.0000000000000142 =  1 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = 0+1i 
assign Y[4'b0100] [46] = 146'h 0000000000000000000000000000040000000;  // +0.0000000000000071 =  1 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = 0+1i 
assign Y[4'b0100] [47] = 146'h 0000000000000000000000000000010000000;  // +0.0000000000000036 =  1 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = 0+1i 
assign Y[4'b0100] [48] = 146'h 0000000000000000000000000000004000000;  // +0.0000000000000018 =  1 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = 0+1i 
assign Y[4'b0100] [49] = 146'h 0000000000000000000000000000001000000;  // +0.0000000000000009 =  1 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = 0+1i 
assign Y[4'b0100] [50] = 146'h 0000000000000000000000000000000400000;  // +0.0000000000000004 =  1 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = 0+1i 
assign Y[4'b0100] [51] = 146'h 0000000000000000000000000000000100000;  // +0.0000000000000002 =  1 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = 0+1i 
assign Y[4'b0100] [52] = 146'h 0000000000000000000000000000000040000;  // +0.0000000000000001 =  1 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = 0+1i 
assign Y[4'b0100] [53] = 146'h 0000000000000000000000000000000010000;  // +0.0000000000000001 =  1 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = 0+1i 
assign Y[4'b0100] [54] = 146'h 0000000000000000000000000000000004000;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = 0+1i 
assign Y[4'b0100] [55] = 146'h 0000000000000000000000000000000001000;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = 0+1i 
assign Y[4'b0100] [56] = 146'h 0000000000000000000000000000000000400;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = 0+1i 
assign Y[4'b0100] [57] = 146'h 0000000000000000000000000000000000100;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = 0+1i 
assign Y[4'b0100] [58] = 146'h 0000000000000000000000000000000000040;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = 0+1i 
assign Y[4'b0100] [59] = 146'h 0000000000000000000000000000000000010;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = 0+1i 
assign Y[4'b0100] [60] = 146'h 0000000000000000000000000000000000004;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = 0+1i 
assign Y[4'b0100] [61] = 146'h 0000000000000000000000000000000000001;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = 0+1i 
assign Y[4'b0100] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = 0+1i 
assign Y[4'b0100] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = 0+1i 
assign Y[4'b0101] [00] = 146'h 00000011044C0C100C4100000000000000000;  // +0.3217505543966422 =  1 * atan( 1 / (  1 + 2^1 ) )   n =  1   d_n = 1+1i 
assign Y[4'b0101] [01] = 146'h 0000001304404040100300000000000000000;  // +0.1973955598498807 =  1 * atan( 1 / (  1 + 2^2 ) )   n =  2   d_n = 1+1i 
assign Y[4'b0101] [02] = 146'h 00000004301110004004C0000000000000000;  // +0.1106572211738956 =  1 * atan( 1 / (  1 + 2^3 ) )   n =  3   d_n = 1+1i 
assign Y[4'b0101] [03] = 146'h 0000000103004444030400000000000000000;  // +0.0587558227157227 =  1 * atan( 1 / (  1 + 2^4 ) )   n =  4   d_n = 1+1i 
assign Y[4'b0101] [04] = 146'h 0000000040300111110310000000000000000;  // +0.0302937599187751 =  1 * atan( 1 / (  1 + 2^5 ) )   n =  5   d_n = 1+1i 
assign Y[4'b0101] [05] = 146'h 0000000010030004444441000000000000000;  // +0.0153834017805952 =  1 * atan( 1 / (  1 + 2^6 ) )   n =  6   d_n = 1+1i 
assign Y[4'b0101] [06] = 146'h 0000000004003000111111000000000000000;  // +0.0077517827122069 =  1 * atan( 1 / (  1 + 2^7 ) )   n =  7   d_n = 1+1i 
assign Y[4'b0101] [07] = 146'h 0000000001000300004444400000000000000;  // +0.0038910309466445 =  1 * atan( 1 / (  1 + 2^8 ) )   n =  8   d_n = 1+1i 
assign Y[4'b0101] [08] = 146'h 0000000000400030000111100000000000000;  // +0.0019493152697654 =  1 * atan( 1 / (  1 + 2^9 ) )   n =  9   d_n = 1+1i 
assign Y[4'b0101] [09] = 146'h 0000000000100003000004440000000000000;  // +0.0009756094465646 =  1 * atan( 1 / (  1 + 2^10 ) )   n = 10   d_n = 1+1i 
assign Y[4'b0101] [10] = 146'h 0000000000040000300000110000000000000;  // +0.0004880429090311 =  1 * atan( 1 / (  1 + 2^11 ) )   n = 11   d_n = 1+1i 
assign Y[4'b0101] [11] = 146'h 0000000000010000030000004000000000000;  // +0.0002440810300565 =  1 * atan( 1 / (  1 + 2^12 ) )   n = 12   d_n = 1+1i 
assign Y[4'b0101] [12] = 146'h 0000000000004000003000000000000000000;  // +0.0001220554125515 =  1 * atan( 1 / (  1 + 2^13 ) )   n = 13   d_n = 1+1i 
assign Y[4'b0101] [13] = 146'h 0000000000001000000300000000000000000;  // +0.0000610314311113 =  1 * atan( 1 / (  1 + 2^14 ) )   n = 14   d_n = 1+1i 
assign Y[4'b0101] [14] = 146'h 0000000000000400000030000000000000000;  // +0.0000305166468214 =  1 * atan( 1 / (  1 + 2^15 ) )   n = 15   d_n = 1+1i 
assign Y[4'b0101] [15] = 146'h 0000000000000100000003000000000000000;  // +0.0000152585562342 =  1 * atan( 1 / (  1 + 2^16 ) )   n = 16   d_n = 1+1i 
assign Y[4'b0101] [16] = 146'h 0000000000000040000000300000000000000;  // +0.0000076293363239 =  1 * atan( 1 / (  1 + 2^17 ) )   n = 17   d_n = 1+1i 
assign Y[4'b0101] [17] = 146'h 0000000000000010000000030000000000000;  // +0.0000038146827137 =  1 * atan( 1 / (  1 + 2^18 ) )   n = 18   d_n = 1+1i 
assign Y[4'b0101] [18] = 146'h 0000000000000004000000003000000000000;  // +0.0000019073449948 =  1 * atan( 1 / (  1 + 2^19 ) )   n = 19   d_n = 1+1i 
assign Y[4'b0101] [19] = 146'h 0000000000000001000000000300000000000;  // +0.0000009536734069 =  1 * atan( 1 / (  1 + 2^20 ) )   n = 20   d_n = 1+1i 
assign Y[4'b0101] [20] = 146'h 0000000000000000400000000030000000000;  // +0.0000004768369308 =  1 * atan( 1 / (  1 + 2^21 ) )   n = 21   d_n = 1+1i 
assign Y[4'b0101] [21] = 146'h 0000000000000000100000000003000000000;  // +0.0000002384185223 =  1 * atan( 1 / (  1 + 2^22 ) )   n = 22   d_n = 1+1i 
assign Y[4'b0101] [22] = 146'h 0000000000000000040000000000300000000;  // +0.0000001192092753 =  1 * atan( 1 / (  1 + 2^23 ) )   n = 23   d_n = 1+1i 
assign Y[4'b0101] [23] = 146'h 0000000000000000010000000000030000000;  // +0.0000000596046412 =  1 * atan( 1 / (  1 + 2^24 ) )   n = 24   d_n = 1+1i 
assign Y[4'b0101] [24] = 146'h 0000000000000000004000000000003000000;  // +0.0000000298023215 =  1 * atan( 1 / (  1 + 2^25 ) )   n = 25   d_n = 1+1i 
assign Y[4'b0101] [25] = 146'h 0000000000000000001000000000000300000;  // +0.0000000149011610 =  1 * atan( 1 / (  1 + 2^26 ) )   n = 26   d_n = 1+1i 
assign Y[4'b0101] [26] = 146'h 0000000000000000000400000000000040000;  // +0.0000000074505805 =  1 * atan( 1 / (  1 + 2^27 ) )   n = 27   d_n = 1+1i 
assign Y[4'b0101] [27] = 146'h 0000000000000000000100000000000000000;  // +0.0000000037252903 =  1 * atan( 1 / (  1 + 2^28 ) )   n = 28   d_n = 1+1i 
assign Y[4'b0101] [28] = 146'h 0000000000000000000040000000000000000;  // +0.0000000018626451 =  1 * atan( 1 / (  1 + 2^29 ) )   n = 29   d_n = 1+1i 
assign Y[4'b0101] [29] = 146'h 0000000000000000000010000000000000000;  // +0.0000000009313226 =  1 * atan( 1 / (  1 + 2^30 ) )   n = 30   d_n = 1+1i 
assign Y[4'b0101] [30] = 146'h 0000000000000000000004000000000000000;  // +0.0000000004656613 =  1 * atan( 1 / (  1 + 2^31 ) )   n = 31   d_n = 1+1i 
assign Y[4'b0101] [31] = 146'h 0000000000000000000001000000000000000;  // +0.0000000002328306 =  1 * atan( 1 / (  1 + 2^32 ) )   n = 32   d_n = 1+1i 
assign Y[4'b0101] [32] = 146'h 0000000000000000000000400000000000000;  // +0.0000000001164153 =  1 * atan( 1 / (  1 + 2^33 ) )   n = 33   d_n = 1+1i 
assign Y[4'b0101] [33] = 146'h 0000000000000000000000100000000000000;  // +0.0000000000582077 =  1 * atan( 1 / (  1 + 2^34 ) )   n = 34   d_n = 1+1i 
assign Y[4'b0101] [34] = 146'h 0000000000000000000000040000000000000;  // +0.0000000000291038 =  1 * atan( 1 / (  1 + 2^35 ) )   n = 35   d_n = 1+1i 
assign Y[4'b0101] [35] = 146'h 0000000000000000000000010000000000000;  // +0.0000000000145519 =  1 * atan( 1 / (  1 + 2^36 ) )   n = 36   d_n = 1+1i 
assign Y[4'b0101] [36] = 146'h 0000000000000000000000004000000000000;  // +0.0000000000072760 =  1 * atan( 1 / (  1 + 2^37 ) )   n = 37   d_n = 1+1i 
assign Y[4'b0101] [37] = 146'h 0000000000000000000000001000000000000;  // +0.0000000000036380 =  1 * atan( 1 / (  1 + 2^38 ) )   n = 38   d_n = 1+1i 
assign Y[4'b0101] [38] = 146'h 0000000000000000000000000400000000000;  // +0.0000000000018190 =  1 * atan( 1 / (  1 + 2^39 ) )   n = 39   d_n = 1+1i 
assign Y[4'b0101] [39] = 146'h 0000000000000000000000000100000000000;  // +0.0000000000009095 =  1 * atan( 1 / (  1 + 2^40 ) )   n = 40   d_n = 1+1i 
assign Y[4'b0101] [40] = 146'h 0000000000000000000000000040000000000;  // +0.0000000000004547 =  1 * atan( 1 / (  1 + 2^41 ) )   n = 41   d_n = 1+1i 
assign Y[4'b0101] [41] = 146'h 0000000000000000000000000010000000000;  // +0.0000000000002274 =  1 * atan( 1 / (  1 + 2^42 ) )   n = 42   d_n = 1+1i 
assign Y[4'b0101] [42] = 146'h 0000000000000000000000000004000000000;  // +0.0000000000001137 =  1 * atan( 1 / (  1 + 2^43 ) )   n = 43   d_n = 1+1i 
assign Y[4'b0101] [43] = 146'h 0000000000000000000000000001000000000;  // +0.0000000000000568 =  1 * atan( 1 / (  1 + 2^44 ) )   n = 44   d_n = 1+1i 
assign Y[4'b0101] [44] = 146'h 0000000000000000000000000000400000000;  // +0.0000000000000284 =  1 * atan( 1 / (  1 + 2^45 ) )   n = 45   d_n = 1+1i 
assign Y[4'b0101] [45] = 146'h 0000000000000000000000000000100000000;  // +0.0000000000000142 =  1 * atan( 1 / (  1 + 2^46 ) )   n = 46   d_n = 1+1i 
assign Y[4'b0101] [46] = 146'h 0000000000000000000000000000040000000;  // +0.0000000000000071 =  1 * atan( 1 / (  1 + 2^47 ) )   n = 47   d_n = 1+1i 
assign Y[4'b0101] [47] = 146'h 0000000000000000000000000000010000000;  // +0.0000000000000036 =  1 * atan( 1 / (  1 + 2^48 ) )   n = 48   d_n = 1+1i 
assign Y[4'b0101] [48] = 146'h 0000000000000000000000000000004000000;  // +0.0000000000000018 =  1 * atan( 1 / (  1 + 2^49 ) )   n = 49   d_n = 1+1i 
assign Y[4'b0101] [49] = 146'h 0000000000000000000000000000001000000;  // +0.0000000000000009 =  1 * atan( 1 / (  1 + 2^50 ) )   n = 50   d_n = 1+1i 
assign Y[4'b0101] [50] = 146'h 0000000000000000000000000000000400000;  // +0.0000000000000004 =  1 * atan( 1 / (  1 + 2^51 ) )   n = 51   d_n = 1+1i 
assign Y[4'b0101] [51] = 146'h 0000000000000000000000000000000100000;  // +0.0000000000000002 =  1 * atan( 1 / (  1 + 2^52 ) )   n = 52   d_n = 1+1i 
assign Y[4'b0101] [52] = 146'h 0000000000000000000000000000000040000;  // +0.0000000000000001 =  1 * atan( 1 / (  1 + 2^53 ) )   n = 53   d_n = 1+1i 
assign Y[4'b0101] [53] = 146'h 0000000000000000000000000000000010000;  // +0.0000000000000001 =  1 * atan( 1 / (  1 + 2^54 ) )   n = 54   d_n = 1+1i 
assign Y[4'b0101] [54] = 146'h 0000000000000000000000000000000004000;  // +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^55 ) )   n = 55   d_n = 1+1i 
assign Y[4'b0101] [55] = 146'h 0000000000000000000000000000000001000;  // +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^56 ) )   n = 56   d_n = 1+1i 
assign Y[4'b0101] [56] = 146'h 0000000000000000000000000000000000400;  // +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^57 ) )   n = 57   d_n = 1+1i 
assign Y[4'b0101] [57] = 146'h 0000000000000000000000000000000000100;  // +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^58 ) )   n = 58   d_n = 1+1i 
assign Y[4'b0101] [58] = 146'h 0000000000000000000000000000000000040;  // +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^59 ) )   n = 59   d_n = 1+1i 
assign Y[4'b0101] [59] = 146'h 0000000000000000000000000000000000010;  // +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^60 ) )   n = 60   d_n = 1+1i 
assign Y[4'b0101] [60] = 146'h 0000000000000000000000000000000000004;  // +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^61 ) )   n = 61   d_n = 1+1i 
assign Y[4'b0101] [61] = 146'h 0000000000000000000000000000000000001;  // +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^62 ) )   n = 62   d_n = 1+1i 
assign Y[4'b0101] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^63 ) )   n = 63   d_n = 1+1i 
assign Y[4'b0101] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^64 ) )   n = 64   d_n = 1+1i 
assign Y[4'b0110] [00] = 146'h 00000040C33304C4300400000000000000000;  // +0.4636476090008061 =  1 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = 0+1i 
assign Y[4'b0110] [01] = 146'h 000000100330C303300300000000000000000;  // +0.2449786631268641 =  1 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = 0+1i 
assign Y[4'b0110] [02] = 146'h 00000004000CCC30C44440000000000000000;  // +0.1243549945467614 =  1 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = 0+1i 
assign Y[4'b0110] [03] = 146'h 00000001000033330C0C30000000000000000;  // +0.0624188099959574 =  1 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = 0+1i 
assign Y[4'b0110] [04] = 146'h 00000000400000CCCCC304000000000000000;  // +0.0312398334302683 =  1 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = 0+1i 
assign Y[4'b0110] [05] = 146'h 0000000010000003333331000000000000000;  // +0.0156237286204768 =  1 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = 0+1i 
assign Y[4'b0110] [06] = 146'h 00000000040000000CCCCCC00000000000000;  // +0.0078123410601011 =  1 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = 0+1i 
assign Y[4'b0110] [07] = 146'h 0000000001000000003333300000000000000;  // +0.0039062301319670 =  1 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = 0+1i 
assign Y[4'b0110] [08] = 146'h 00000000004000000000CCCC0000000000000;  // +0.0019531225164788 =  1 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = 0+1i 
assign Y[4'b0110] [09] = 146'h 0000000000100000000003330000000000000;  // +0.0009765621895593 =  1 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = 0+1i 
assign Y[4'b0110] [10] = 146'h 00000000000400000000000CC000000000000;  // +0.0004882812111949 =  1 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = 0+1i 
assign Y[4'b0110] [11] = 146'h 0000000000010000000000003000000000000;  // +0.0002441406201494 =  1 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = 0+1i 
assign Y[4'b0110] [12] = 146'h 0000000000004000000000000400000000000;  // +0.0001220703118937 =  1 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = 0+1i 
assign Y[4'b0110] [13] = 146'h 0000000000001000000000000000000000000;  // +0.0000610351561742 =  1 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = 0+1i 
assign Y[4'b0110] [14] = 146'h 0000000000000400000000000000000000000;  // +0.0000305175781155 =  1 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = 0+1i 
assign Y[4'b0110] [15] = 146'h 0000000000000100000000000000000000000;  // +0.0000152587890613 =  1 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = 0+1i 
assign Y[4'b0110] [16] = 146'h 0000000000000040000000000000000000000;  // +0.0000076293945311 =  1 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = 0+1i 
assign Y[4'b0110] [17] = 146'h 0000000000000010000000000000000000000;  // +0.0000038146972656 =  1 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = 0+1i 
assign Y[4'b0110] [18] = 146'h 0000000000000004000000000000000000000;  // +0.0000019073486328 =  1 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = 0+1i 
assign Y[4'b0110] [19] = 146'h 0000000000000001000000000000000000000;  // +0.0000009536743164 =  1 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = 0+1i 
assign Y[4'b0110] [20] = 146'h 0000000000000000400000000000000000000;  // +0.0000004768371582 =  1 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = 0+1i 
assign Y[4'b0110] [21] = 146'h 0000000000000000100000000000000000000;  // +0.0000002384185791 =  1 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = 0+1i 
assign Y[4'b0110] [22] = 146'h 0000000000000000040000000000000000000;  // +0.0000001192092896 =  1 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = 0+1i 
assign Y[4'b0110] [23] = 146'h 0000000000000000010000000000000000000;  // +0.0000000596046448 =  1 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = 0+1i 
assign Y[4'b0110] [24] = 146'h 0000000000000000004000000000000000000;  // +0.0000000298023224 =  1 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = 0+1i 
assign Y[4'b0110] [25] = 146'h 0000000000000000001000000000000000000;  // +0.0000000149011612 =  1 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = 0+1i 
assign Y[4'b0110] [26] = 146'h 0000000000000000000400000000000000000;  // +0.0000000074505806 =  1 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = 0+1i 
assign Y[4'b0110] [27] = 146'h 0000000000000000000100000000000000000;  // +0.0000000037252903 =  1 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = 0+1i 
assign Y[4'b0110] [28] = 146'h 0000000000000000000040000000000000000;  // +0.0000000018626451 =  1 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = 0+1i 
assign Y[4'b0110] [29] = 146'h 0000000000000000000010000000000000000;  // +0.0000000009313226 =  1 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = 0+1i 
assign Y[4'b0110] [30] = 146'h 0000000000000000000004000000000000000;  // +0.0000000004656613 =  1 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = 0+1i 
assign Y[4'b0110] [31] = 146'h 0000000000000000000001000000000000000;  // +0.0000000002328306 =  1 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = 0+1i 
assign Y[4'b0110] [32] = 146'h 0000000000000000000000400000000000000;  // +0.0000000001164153 =  1 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = 0+1i 
assign Y[4'b0110] [33] = 146'h 0000000000000000000000100000000000000;  // +0.0000000000582077 =  1 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = 0+1i 
assign Y[4'b0110] [34] = 146'h 0000000000000000000000040000000000000;  // +0.0000000000291038 =  1 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = 0+1i 
assign Y[4'b0110] [35] = 146'h 0000000000000000000000010000000000000;  // +0.0000000000145519 =  1 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = 0+1i 
assign Y[4'b0110] [36] = 146'h 0000000000000000000000004000000000000;  // +0.0000000000072760 =  1 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = 0+1i 
assign Y[4'b0110] [37] = 146'h 0000000000000000000000001000000000000;  // +0.0000000000036380 =  1 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = 0+1i 
assign Y[4'b0110] [38] = 146'h 0000000000000000000000000400000000000;  // +0.0000000000018190 =  1 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = 0+1i 
assign Y[4'b0110] [39] = 146'h 0000000000000000000000000100000000000;  // +0.0000000000009095 =  1 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = 0+1i 
assign Y[4'b0110] [40] = 146'h 0000000000000000000000000040000000000;  // +0.0000000000004547 =  1 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = 0+1i 
assign Y[4'b0110] [41] = 146'h 0000000000000000000000000010000000000;  // +0.0000000000002274 =  1 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = 0+1i 
assign Y[4'b0110] [42] = 146'h 0000000000000000000000000004000000000;  // +0.0000000000001137 =  1 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = 0+1i 
assign Y[4'b0110] [43] = 146'h 0000000000000000000000000001000000000;  // +0.0000000000000568 =  1 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = 0+1i 
assign Y[4'b0110] [44] = 146'h 0000000000000000000000000000400000000;  // +0.0000000000000284 =  1 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = 0+1i 
assign Y[4'b0110] [45] = 146'h 0000000000000000000000000000100000000;  // +0.0000000000000142 =  1 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = 0+1i 
assign Y[4'b0110] [46] = 146'h 0000000000000000000000000000040000000;  // +0.0000000000000071 =  1 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = 0+1i 
assign Y[4'b0110] [47] = 146'h 0000000000000000000000000000010000000;  // +0.0000000000000036 =  1 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = 0+1i 
assign Y[4'b0110] [48] = 146'h 0000000000000000000000000000004000000;  // +0.0000000000000018 =  1 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = 0+1i 
assign Y[4'b0110] [49] = 146'h 0000000000000000000000000000001000000;  // +0.0000000000000009 =  1 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = 0+1i 
assign Y[4'b0110] [50] = 146'h 0000000000000000000000000000000400000;  // +0.0000000000000004 =  1 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = 0+1i 
assign Y[4'b0110] [51] = 146'h 0000000000000000000000000000000100000;  // +0.0000000000000002 =  1 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = 0+1i 
assign Y[4'b0110] [52] = 146'h 0000000000000000000000000000000040000;  // +0.0000000000000001 =  1 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = 0+1i 
assign Y[4'b0110] [53] = 146'h 0000000000000000000000000000000010000;  // +0.0000000000000001 =  1 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = 0+1i 
assign Y[4'b0110] [54] = 146'h 0000000000000000000000000000000004000;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = 0+1i 
assign Y[4'b0110] [55] = 146'h 0000000000000000000000000000000001000;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = 0+1i 
assign Y[4'b0110] [56] = 146'h 0000000000000000000000000000000000400;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = 0+1i 
assign Y[4'b0110] [57] = 146'h 0000000000000000000000000000000000100;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = 0+1i 
assign Y[4'b0110] [58] = 146'h 0000000000000000000000000000000000040;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = 0+1i 
assign Y[4'b0110] [59] = 146'h 0000000000000000000000000000000000010;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = 0+1i 
assign Y[4'b0110] [60] = 146'h 0000000000000000000000000000000000004;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = 0+1i 
assign Y[4'b0110] [61] = 146'h 0000000000000000000000000000000000001;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = 0+1i 
assign Y[4'b0110] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = 0+1i 
assign Y[4'b0110] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = 0+1i 
assign Y[4'b0111] [00] = 146'h 000001304101000CC44000000000000000000;  // +0.7853981633974483 =  1 * atan( 1 / ( -1 + 2^1 ) )   n =  1   d_n = -1+1i 
assign Y[4'b0111] [01] = 146'h 00000011044C0C100C4100000000000000000;  // +0.3217505543966422 =  1 * atan( 1 / ( -1 + 2^2 ) )   n =  2   d_n = -1+1i 
assign Y[4'b0111] [02] = 146'h 00000004101110CC0CC040000000000000000;  // +0.1418970546041639 =  1 * atan( 1 / ( -1 + 2^3 ) )   n =  3   d_n = -1+1i 
assign Y[4'b0111] [03] = 146'h 00000001010044443040D0000000000000000;  // +0.0665681637758238 =  1 * atan( 1 / ( -1 + 2^4 ) )   n =  4   d_n = -1+1i 
assign Y[4'b0111] [04] = 146'h 0000000040100111110C44000000000000000;  // +0.0322468824352539 =  1 * atan( 1 / ( -1 + 2^5 ) )   n =  5   d_n = -1+1i 
assign Y[4'b0111] [05] = 146'h 0000000010010004444441000000000000000;  // +0.0158716829917901 =  1 * atan( 1 / ( -1 + 2^6 ) )   n =  6   d_n = -1+1i 
assign Y[4'b0111] [06] = 146'h 0000000004001000111111000000000000000;  // +0.0078738530241005 =  1 * atan( 1 / ( -1 + 2^7 ) )   n =  7   d_n = -1+1i 
assign Y[4'b0111] [07] = 146'h 0000000001000100004444400000000000000;  // +0.0039215485247600 =  1 * atan( 1 / ( -1 + 2^8 ) )   n =  8   d_n = -1+1i 
assign Y[4'b0111] [08] = 146'h 0000000000400010000111100000000000000;  // +0.0019569446642965 =  1 * atan( 1 / ( -1 + 2^9 ) )   n =  9   d_n = -1+1i 
assign Y[4'b0111] [09] = 146'h 0000000000100001000004440000000000000;  // +0.0009775167951974 =  1 * atan( 1 / ( -1 + 2^10 ) )   n = 10   d_n = -1+1i 
assign Y[4'b0111] [10] = 146'h 0000000000040000100000110000000000000;  // +0.0004885197461893 =  1 * atan( 1 / ( -1 + 2^11 ) )   n = 11   d_n = -1+1i 
assign Y[4'b0111] [11] = 146'h 0000000000010000010000004000000000000;  // +0.0002442002393461 =  1 * atan( 1 / ( -1 + 2^12 ) )   n = 12   d_n = -1+1i 
assign Y[4'b0111] [12] = 146'h 0000000000004000001000000000000000000;  // +0.0001220852148739 =  1 * atan( 1 / ( -1 + 2^13 ) )   n = 13   d_n = -1+1i 
assign Y[4'b0111] [13] = 146'h 0000000000001000000100000000000000000;  // +0.0000610388816919 =  1 * atan( 1 / ( -1 + 2^14 ) )   n = 14   d_n = -1+1i 
assign Y[4'b0111] [14] = 146'h 0000000000000400000010000000000000000;  // +0.0000305185094665 =  1 * atan( 1 / ( -1 + 2^15 ) )   n = 15   d_n = -1+1i 
assign Y[4'b0111] [15] = 146'h 0000000000000100000001000000000000000;  // +0.0000152590218955 =  1 * atan( 1 / ( -1 + 2^16 ) )   n = 16   d_n = -1+1i 
assign Y[4'b0111] [16] = 146'h 0000000000000040000000100000000000000;  // +0.0000076294527392 =  1 * atan( 1 / ( -1 + 2^17 ) )   n = 17   d_n = -1+1i 
assign Y[4'b0111] [17] = 146'h 0000000000000010000000010000000000000;  // +0.0000038147118176 =  1 * atan( 1 / ( -1 + 2^18 ) )   n = 18   d_n = -1+1i 
assign Y[4'b0111] [18] = 146'h 0000000000000004000000001000000000000;  // +0.0000019073522708 =  1 * atan( 1 / ( -1 + 2^19 ) )   n = 19   d_n = -1+1i 
assign Y[4'b0111] [19] = 146'h 0000000000000001000000000100000000000;  // +0.0000009536752259 =  1 * atan( 1 / ( -1 + 2^20 ) )   n = 20   d_n = -1+1i 
assign Y[4'b0111] [20] = 146'h 0000000000000000400000000010000000000;  // +0.0000004768373856 =  1 * atan( 1 / ( -1 + 2^21 ) )   n = 21   d_n = -1+1i 
assign Y[4'b0111] [21] = 146'h 0000000000000000100000000001000000000;  // +0.0000002384186359 =  1 * atan( 1 / ( -1 + 2^22 ) )   n = 22   d_n = -1+1i 
assign Y[4'b0111] [22] = 146'h 0000000000000000040000000000100000000;  // +0.0000001192093038 =  1 * atan( 1 / ( -1 + 2^23 ) )   n = 23   d_n = -1+1i 
assign Y[4'b0111] [23] = 146'h 0000000000000000010000000000010000000;  // +0.0000000596046483 =  1 * atan( 1 / ( -1 + 2^24 ) )   n = 24   d_n = -1+1i 
assign Y[4'b0111] [24] = 146'h 0000000000000000004000000000001000000;  // +0.0000000298023233 =  1 * atan( 1 / ( -1 + 2^25 ) )   n = 25   d_n = -1+1i 
assign Y[4'b0111] [25] = 146'h 0000000000000000001000000000000100000;  // +0.0000000149011614 =  1 * atan( 1 / ( -1 + 2^26 ) )   n = 26   d_n = -1+1i 
assign Y[4'b0111] [26] = 146'h 0000000000000000000400000000000000000;  // +0.0000000074505807 =  1 * atan( 1 / ( -1 + 2^27 ) )   n = 27   d_n = -1+1i 
assign Y[4'b0111] [27] = 146'h 0000000000000000000100000000000000000;  // +0.0000000037252903 =  1 * atan( 1 / ( -1 + 2^28 ) )   n = 28   d_n = -1+1i 
assign Y[4'b0111] [28] = 146'h 0000000000000000000040000000000000000;  // +0.0000000018626452 =  1 * atan( 1 / ( -1 + 2^29 ) )   n = 29   d_n = -1+1i 
assign Y[4'b0111] [29] = 146'h 0000000000000000000010000000000000000;  // +0.0000000009313226 =  1 * atan( 1 / ( -1 + 2^30 ) )   n = 30   d_n = -1+1i 
assign Y[4'b0111] [30] = 146'h 0000000000000000000004000000000000000;  // +0.0000000004656613 =  1 * atan( 1 / ( -1 + 2^31 ) )   n = 31   d_n = -1+1i 
assign Y[4'b0111] [31] = 146'h 0000000000000000000001000000000000000;  // +0.0000000002328306 =  1 * atan( 1 / ( -1 + 2^32 ) )   n = 32   d_n = -1+1i 
assign Y[4'b0111] [32] = 146'h 0000000000000000000000400000000000000;  // +0.0000000001164153 =  1 * atan( 1 / ( -1 + 2^33 ) )   n = 33   d_n = -1+1i 
assign Y[4'b0111] [33] = 146'h 0000000000000000000000100000000000000;  // +0.0000000000582077 =  1 * atan( 1 / ( -1 + 2^34 ) )   n = 34   d_n = -1+1i 
assign Y[4'b0111] [34] = 146'h 0000000000000000000000040000000000000;  // +0.0000000000291038 =  1 * atan( 1 / ( -1 + 2^35 ) )   n = 35   d_n = -1+1i 
assign Y[4'b0111] [35] = 146'h 0000000000000000000000010000000000000;  // +0.0000000000145519 =  1 * atan( 1 / ( -1 + 2^36 ) )   n = 36   d_n = -1+1i 
assign Y[4'b0111] [36] = 146'h 0000000000000000000000004000000000000;  // +0.0000000000072760 =  1 * atan( 1 / ( -1 + 2^37 ) )   n = 37   d_n = -1+1i 
assign Y[4'b0111] [37] = 146'h 0000000000000000000000001000000000000;  // +0.0000000000036380 =  1 * atan( 1 / ( -1 + 2^38 ) )   n = 38   d_n = -1+1i 
assign Y[4'b0111] [38] = 146'h 0000000000000000000000000400000000000;  // +0.0000000000018190 =  1 * atan( 1 / ( -1 + 2^39 ) )   n = 39   d_n = -1+1i 
assign Y[4'b0111] [39] = 146'h 0000000000000000000000000100000000000;  // +0.0000000000009095 =  1 * atan( 1 / ( -1 + 2^40 ) )   n = 40   d_n = -1+1i 
assign Y[4'b0111] [40] = 146'h 0000000000000000000000000040000000000;  // +0.0000000000004547 =  1 * atan( 1 / ( -1 + 2^41 ) )   n = 41   d_n = -1+1i 
assign Y[4'b0111] [41] = 146'h 0000000000000000000000000010000000000;  // +0.0000000000002274 =  1 * atan( 1 / ( -1 + 2^42 ) )   n = 42   d_n = -1+1i 
assign Y[4'b0111] [42] = 146'h 0000000000000000000000000004000000000;  // +0.0000000000001137 =  1 * atan( 1 / ( -1 + 2^43 ) )   n = 43   d_n = -1+1i 
assign Y[4'b0111] [43] = 146'h 0000000000000000000000000001000000000;  // +0.0000000000000568 =  1 * atan( 1 / ( -1 + 2^44 ) )   n = 44   d_n = -1+1i 
assign Y[4'b0111] [44] = 146'h 0000000000000000000000000000400000000;  // +0.0000000000000284 =  1 * atan( 1 / ( -1 + 2^45 ) )   n = 45   d_n = -1+1i 
assign Y[4'b0111] [45] = 146'h 0000000000000000000000000000100000000;  // +0.0000000000000142 =  1 * atan( 1 / ( -1 + 2^46 ) )   n = 46   d_n = -1+1i 
assign Y[4'b0111] [46] = 146'h 0000000000000000000000000000040000000;  // +0.0000000000000071 =  1 * atan( 1 / ( -1 + 2^47 ) )   n = 47   d_n = -1+1i 
assign Y[4'b0111] [47] = 146'h 0000000000000000000000000000010000000;  // +0.0000000000000036 =  1 * atan( 1 / ( -1 + 2^48 ) )   n = 48   d_n = -1+1i 
assign Y[4'b0111] [48] = 146'h 0000000000000000000000000000004000000;  // +0.0000000000000018 =  1 * atan( 1 / ( -1 + 2^49 ) )   n = 49   d_n = -1+1i 
assign Y[4'b0111] [49] = 146'h 0000000000000000000000000000001000000;  // +0.0000000000000009 =  1 * atan( 1 / ( -1 + 2^50 ) )   n = 50   d_n = -1+1i 
assign Y[4'b0111] [50] = 146'h 0000000000000000000000000000000400000;  // +0.0000000000000004 =  1 * atan( 1 / ( -1 + 2^51 ) )   n = 51   d_n = -1+1i 
assign Y[4'b0111] [51] = 146'h 0000000000000000000000000000000100000;  // +0.0000000000000002 =  1 * atan( 1 / ( -1 + 2^52 ) )   n = 52   d_n = -1+1i 
assign Y[4'b0111] [52] = 146'h 0000000000000000000000000000000040000;  // +0.0000000000000001 =  1 * atan( 1 / ( -1 + 2^53 ) )   n = 53   d_n = -1+1i 
assign Y[4'b0111] [53] = 146'h 0000000000000000000000000000000010000;  // +0.0000000000000001 =  1 * atan( 1 / ( -1 + 2^54 ) )   n = 54   d_n = -1+1i 
assign Y[4'b0111] [54] = 146'h 0000000000000000000000000000000004000;  // +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^55 ) )   n = 55   d_n = -1+1i 
assign Y[4'b0111] [55] = 146'h 0000000000000000000000000000000001000;  // +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^56 ) )   n = 56   d_n = -1+1i 
assign Y[4'b0111] [56] = 146'h 0000000000000000000000000000000000400;  // +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^57 ) )   n = 57   d_n = -1+1i 
assign Y[4'b0111] [57] = 146'h 0000000000000000000000000000000000100;  // +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^58 ) )   n = 58   d_n = -1+1i 
assign Y[4'b0111] [58] = 146'h 0000000000000000000000000000000000040;  // +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^59 ) )   n = 59   d_n = -1+1i 
assign Y[4'b0111] [59] = 146'h 0000000000000000000000000000000000010;  // +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^60 ) )   n = 60   d_n = -1+1i 
assign Y[4'b0111] [60] = 146'h 0000000000000000000000000000000000004;  // +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^61 ) )   n = 61   d_n = -1+1i 
assign Y[4'b0111] [61] = 146'h 0000000000000000000000000000000000001;  // +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^62 ) )   n = 62   d_n = -1+1i 
assign Y[4'b0111] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^63 ) )   n = 63   d_n = -1+1i 
assign Y[4'b0111] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^64 ) )   n = 64   d_n = -1+1i 
assign Y[4'b1000] [00] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = 0 
assign Y[4'b1000] [01] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = 0 
assign Y[4'b1000] [02] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = 0 
assign Y[4'b1000] [03] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = 0 
assign Y[4'b1000] [04] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = 0 
assign Y[4'b1000] [05] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = 0 
assign Y[4'b1000] [06] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = 0 
assign Y[4'b1000] [07] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = 0 
assign Y[4'b1000] [08] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = 0 
assign Y[4'b1000] [09] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = 0 
assign Y[4'b1000] [10] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = 0 
assign Y[4'b1000] [11] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = 0 
assign Y[4'b1000] [12] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = 0 
assign Y[4'b1000] [13] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = 0 
assign Y[4'b1000] [14] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = 0 
assign Y[4'b1000] [15] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = 0 
assign Y[4'b1000] [16] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = 0 
assign Y[4'b1000] [17] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = 0 
assign Y[4'b1000] [18] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = 0 
assign Y[4'b1000] [19] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = 0 
assign Y[4'b1000] [20] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = 0 
assign Y[4'b1000] [21] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = 0 
assign Y[4'b1000] [22] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = 0 
assign Y[4'b1000] [23] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = 0 
assign Y[4'b1000] [24] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = 0 
assign Y[4'b1000] [25] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = 0 
assign Y[4'b1000] [26] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = 0 
assign Y[4'b1000] [27] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = 0 
assign Y[4'b1000] [28] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = 0 
assign Y[4'b1000] [29] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = 0 
assign Y[4'b1000] [30] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = 0 
assign Y[4'b1000] [31] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = 0 
assign Y[4'b1000] [32] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = 0 
assign Y[4'b1000] [33] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = 0 
assign Y[4'b1000] [34] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = 0 
assign Y[4'b1000] [35] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = 0 
assign Y[4'b1000] [36] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = 0 
assign Y[4'b1000] [37] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = 0 
assign Y[4'b1000] [38] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = 0 
assign Y[4'b1000] [39] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = 0 
assign Y[4'b1000] [40] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = 0 
assign Y[4'b1000] [41] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = 0 
assign Y[4'b1000] [42] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = 0 
assign Y[4'b1000] [43] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = 0 
assign Y[4'b1000] [44] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = 0 
assign Y[4'b1000] [45] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = 0 
assign Y[4'b1000] [46] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = 0 
assign Y[4'b1000] [47] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = 0 
assign Y[4'b1000] [48] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = 0 
assign Y[4'b1000] [49] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = 0 
assign Y[4'b1000] [50] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = 0 
assign Y[4'b1000] [51] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = 0 
assign Y[4'b1000] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = 0 
assign Y[4'b1000] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = 0 
assign Y[4'b1000] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = 0 
assign Y[4'b1000] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = 0 
assign Y[4'b1000] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = 0 
assign Y[4'b1000] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = 0 
assign Y[4'b1000] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = 0 
assign Y[4'b1000] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = 0 
assign Y[4'b1000] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = 0 
assign Y[4'b1000] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = 0 
assign Y[4'b1000] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = 0 
assign Y[4'b1000] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = 0 
assign Y[4'b1001] [00] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^1 ) )   n =  1   d_n = 1 
assign Y[4'b1001] [01] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^2 ) )   n =  2   d_n = 1 
assign Y[4'b1001] [02] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^3 ) )   n =  3   d_n = 1 
assign Y[4'b1001] [03] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^4 ) )   n =  4   d_n = 1 
assign Y[4'b1001] [04] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^5 ) )   n =  5   d_n = 1 
assign Y[4'b1001] [05] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^6 ) )   n =  6   d_n = 1 
assign Y[4'b1001] [06] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^7 ) )   n =  7   d_n = 1 
assign Y[4'b1001] [07] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^8 ) )   n =  8   d_n = 1 
assign Y[4'b1001] [08] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^9 ) )   n =  9   d_n = 1 
assign Y[4'b1001] [09] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^10 ) )   n = 10   d_n = 1 
assign Y[4'b1001] [10] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^11 ) )   n = 11   d_n = 1 
assign Y[4'b1001] [11] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^12 ) )   n = 12   d_n = 1 
assign Y[4'b1001] [12] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^13 ) )   n = 13   d_n = 1 
assign Y[4'b1001] [13] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^14 ) )   n = 14   d_n = 1 
assign Y[4'b1001] [14] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^15 ) )   n = 15   d_n = 1 
assign Y[4'b1001] [15] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^16 ) )   n = 16   d_n = 1 
assign Y[4'b1001] [16] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^17 ) )   n = 17   d_n = 1 
assign Y[4'b1001] [17] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^18 ) )   n = 18   d_n = 1 
assign Y[4'b1001] [18] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^19 ) )   n = 19   d_n = 1 
assign Y[4'b1001] [19] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^20 ) )   n = 20   d_n = 1 
assign Y[4'b1001] [20] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^21 ) )   n = 21   d_n = 1 
assign Y[4'b1001] [21] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^22 ) )   n = 22   d_n = 1 
assign Y[4'b1001] [22] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^23 ) )   n = 23   d_n = 1 
assign Y[4'b1001] [23] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^24 ) )   n = 24   d_n = 1 
assign Y[4'b1001] [24] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^25 ) )   n = 25   d_n = 1 
assign Y[4'b1001] [25] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^26 ) )   n = 26   d_n = 1 
assign Y[4'b1001] [26] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^27 ) )   n = 27   d_n = 1 
assign Y[4'b1001] [27] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^28 ) )   n = 28   d_n = 1 
assign Y[4'b1001] [28] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^29 ) )   n = 29   d_n = 1 
assign Y[4'b1001] [29] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^30 ) )   n = 30   d_n = 1 
assign Y[4'b1001] [30] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^31 ) )   n = 31   d_n = 1 
assign Y[4'b1001] [31] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^32 ) )   n = 32   d_n = 1 
assign Y[4'b1001] [32] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^33 ) )   n = 33   d_n = 1 
assign Y[4'b1001] [33] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^34 ) )   n = 34   d_n = 1 
assign Y[4'b1001] [34] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^35 ) )   n = 35   d_n = 1 
assign Y[4'b1001] [35] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^36 ) )   n = 36   d_n = 1 
assign Y[4'b1001] [36] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^37 ) )   n = 37   d_n = 1 
assign Y[4'b1001] [37] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^38 ) )   n = 38   d_n = 1 
assign Y[4'b1001] [38] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^39 ) )   n = 39   d_n = 1 
assign Y[4'b1001] [39] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^40 ) )   n = 40   d_n = 1 
assign Y[4'b1001] [40] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^41 ) )   n = 41   d_n = 1 
assign Y[4'b1001] [41] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^42 ) )   n = 42   d_n = 1 
assign Y[4'b1001] [42] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^43 ) )   n = 43   d_n = 1 
assign Y[4'b1001] [43] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^44 ) )   n = 44   d_n = 1 
assign Y[4'b1001] [44] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^45 ) )   n = 45   d_n = 1 
assign Y[4'b1001] [45] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^46 ) )   n = 46   d_n = 1 
assign Y[4'b1001] [46] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^47 ) )   n = 47   d_n = 1 
assign Y[4'b1001] [47] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^48 ) )   n = 48   d_n = 1 
assign Y[4'b1001] [48] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^49 ) )   n = 49   d_n = 1 
assign Y[4'b1001] [49] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^50 ) )   n = 50   d_n = 1 
assign Y[4'b1001] [50] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^51 ) )   n = 51   d_n = 1 
assign Y[4'b1001] [51] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^52 ) )   n = 52   d_n = 1 
assign Y[4'b1001] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^53 ) )   n = 53   d_n = 1 
assign Y[4'b1001] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^54 ) )   n = 54   d_n = 1 
assign Y[4'b1001] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^55 ) )   n = 55   d_n = 1 
assign Y[4'b1001] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^56 ) )   n = 56   d_n = 1 
assign Y[4'b1001] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^57 ) )   n = 57   d_n = 1 
assign Y[4'b1001] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^58 ) )   n = 58   d_n = 1 
assign Y[4'b1001] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^59 ) )   n = 59   d_n = 1 
assign Y[4'b1001] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^60 ) )   n = 60   d_n = 1 
assign Y[4'b1001] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^61 ) )   n = 61   d_n = 1 
assign Y[4'b1001] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^62 ) )   n = 62   d_n = 1 
assign Y[4'b1001] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^63 ) )   n = 63   d_n = 1 
assign Y[4'b1001] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^64 ) )   n = 64   d_n = 1 
assign Y[4'b1010] [00] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = -0 
assign Y[4'b1010] [01] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = -0 
assign Y[4'b1010] [02] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = -0 
assign Y[4'b1010] [03] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = -0 
assign Y[4'b1010] [04] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = -0 
assign Y[4'b1010] [05] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = -0 
assign Y[4'b1010] [06] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = -0 
assign Y[4'b1010] [07] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = -0 
assign Y[4'b1010] [08] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = -0 
assign Y[4'b1010] [09] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = -0 
assign Y[4'b1010] [10] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = -0 
assign Y[4'b1010] [11] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = -0 
assign Y[4'b1010] [12] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = -0 
assign Y[4'b1010] [13] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = -0 
assign Y[4'b1010] [14] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = -0 
assign Y[4'b1010] [15] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = -0 
assign Y[4'b1010] [16] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = -0 
assign Y[4'b1010] [17] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = -0 
assign Y[4'b1010] [18] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = -0 
assign Y[4'b1010] [19] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = -0 
assign Y[4'b1010] [20] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = -0 
assign Y[4'b1010] [21] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = -0 
assign Y[4'b1010] [22] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = -0 
assign Y[4'b1010] [23] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = -0 
assign Y[4'b1010] [24] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = -0 
assign Y[4'b1010] [25] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = -0 
assign Y[4'b1010] [26] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = -0 
assign Y[4'b1010] [27] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = -0 
assign Y[4'b1010] [28] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = -0 
assign Y[4'b1010] [29] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = -0 
assign Y[4'b1010] [30] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = -0 
assign Y[4'b1010] [31] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = -0 
assign Y[4'b1010] [32] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = -0 
assign Y[4'b1010] [33] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = -0 
assign Y[4'b1010] [34] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = -0 
assign Y[4'b1010] [35] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = -0 
assign Y[4'b1010] [36] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = -0 
assign Y[4'b1010] [37] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = -0 
assign Y[4'b1010] [38] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = -0 
assign Y[4'b1010] [39] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = -0 
assign Y[4'b1010] [40] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = -0 
assign Y[4'b1010] [41] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = -0 
assign Y[4'b1010] [42] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = -0 
assign Y[4'b1010] [43] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = -0 
assign Y[4'b1010] [44] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = -0 
assign Y[4'b1010] [45] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = -0 
assign Y[4'b1010] [46] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = -0 
assign Y[4'b1010] [47] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = -0 
assign Y[4'b1010] [48] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = -0 
assign Y[4'b1010] [49] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = -0 
assign Y[4'b1010] [50] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = -0 
assign Y[4'b1010] [51] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = -0 
assign Y[4'b1010] [52] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = -0 
assign Y[4'b1010] [53] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = -0 
assign Y[4'b1010] [54] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = -0 
assign Y[4'b1010] [55] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = -0 
assign Y[4'b1010] [56] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = -0 
assign Y[4'b1010] [57] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = -0 
assign Y[4'b1010] [58] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = -0 
assign Y[4'b1010] [59] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = -0 
assign Y[4'b1010] [60] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = -0 
assign Y[4'b1010] [61] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = -0 
assign Y[4'b1010] [62] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = -0 
assign Y[4'b1010] [63] = 146'h 0000000000000000000000000000000000000;  // +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = -0 
assign Y[4'b1011] [00] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^1 ) )   n =  1   d_n = -1 
assign Y[4'b1011] [01] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^2 ) )   n =  2   d_n = -1 
assign Y[4'b1011] [02] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^3 ) )   n =  3   d_n = -1 
assign Y[4'b1011] [03] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^4 ) )   n =  4   d_n = -1 
assign Y[4'b1011] [04] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^5 ) )   n =  5   d_n = -1 
assign Y[4'b1011] [05] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^6 ) )   n =  6   d_n = -1 
assign Y[4'b1011] [06] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^7 ) )   n =  7   d_n = -1 
assign Y[4'b1011] [07] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^8 ) )   n =  8   d_n = -1 
assign Y[4'b1011] [08] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^9 ) )   n =  9   d_n = -1 
assign Y[4'b1011] [09] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^10 ) )   n = 10   d_n = -1 
assign Y[4'b1011] [10] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^11 ) )   n = 11   d_n = -1 
assign Y[4'b1011] [11] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^12 ) )   n = 12   d_n = -1 
assign Y[4'b1011] [12] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^13 ) )   n = 13   d_n = -1 
assign Y[4'b1011] [13] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^14 ) )   n = 14   d_n = -1 
assign Y[4'b1011] [14] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^15 ) )   n = 15   d_n = -1 
assign Y[4'b1011] [15] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^16 ) )   n = 16   d_n = -1 
assign Y[4'b1011] [16] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^17 ) )   n = 17   d_n = -1 
assign Y[4'b1011] [17] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^18 ) )   n = 18   d_n = -1 
assign Y[4'b1011] [18] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^19 ) )   n = 19   d_n = -1 
assign Y[4'b1011] [19] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^20 ) )   n = 20   d_n = -1 
assign Y[4'b1011] [20] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^21 ) )   n = 21   d_n = -1 
assign Y[4'b1011] [21] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^22 ) )   n = 22   d_n = -1 
assign Y[4'b1011] [22] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^23 ) )   n = 23   d_n = -1 
assign Y[4'b1011] [23] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^24 ) )   n = 24   d_n = -1 
assign Y[4'b1011] [24] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^25 ) )   n = 25   d_n = -1 
assign Y[4'b1011] [25] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^26 ) )   n = 26   d_n = -1 
assign Y[4'b1011] [26] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^27 ) )   n = 27   d_n = -1 
assign Y[4'b1011] [27] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^28 ) )   n = 28   d_n = -1 
assign Y[4'b1011] [28] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^29 ) )   n = 29   d_n = -1 
assign Y[4'b1011] [29] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^30 ) )   n = 30   d_n = -1 
assign Y[4'b1011] [30] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^31 ) )   n = 31   d_n = -1 
assign Y[4'b1011] [31] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^32 ) )   n = 32   d_n = -1 
assign Y[4'b1011] [32] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^33 ) )   n = 33   d_n = -1 
assign Y[4'b1011] [33] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^34 ) )   n = 34   d_n = -1 
assign Y[4'b1011] [34] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^35 ) )   n = 35   d_n = -1 
assign Y[4'b1011] [35] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^36 ) )   n = 36   d_n = -1 
assign Y[4'b1011] [36] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^37 ) )   n = 37   d_n = -1 
assign Y[4'b1011] [37] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^38 ) )   n = 38   d_n = -1 
assign Y[4'b1011] [38] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^39 ) )   n = 39   d_n = -1 
assign Y[4'b1011] [39] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^40 ) )   n = 40   d_n = -1 
assign Y[4'b1011] [40] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^41 ) )   n = 41   d_n = -1 
assign Y[4'b1011] [41] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^42 ) )   n = 42   d_n = -1 
assign Y[4'b1011] [42] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^43 ) )   n = 43   d_n = -1 
assign Y[4'b1011] [43] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^44 ) )   n = 44   d_n = -1 
assign Y[4'b1011] [44] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^45 ) )   n = 45   d_n = -1 
assign Y[4'b1011] [45] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^46 ) )   n = 46   d_n = -1 
assign Y[4'b1011] [46] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^47 ) )   n = 47   d_n = -1 
assign Y[4'b1011] [47] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^48 ) )   n = 48   d_n = -1 
assign Y[4'b1011] [48] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^49 ) )   n = 49   d_n = -1 
assign Y[4'b1011] [49] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^50 ) )   n = 50   d_n = -1 
assign Y[4'b1011] [50] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^51 ) )   n = 51   d_n = -1 
assign Y[4'b1011] [51] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^52 ) )   n = 52   d_n = -1 
assign Y[4'b1011] [52] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^53 ) )   n = 53   d_n = -1 
assign Y[4'b1011] [53] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^54 ) )   n = 54   d_n = -1 
assign Y[4'b1011] [54] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^55 ) )   n = 55   d_n = -1 
assign Y[4'b1011] [55] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^56 ) )   n = 56   d_n = -1 
assign Y[4'b1011] [56] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^57 ) )   n = 57   d_n = -1 
assign Y[4'b1011] [57] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^58 ) )   n = 58   d_n = -1 
assign Y[4'b1011] [58] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^59 ) )   n = 59   d_n = -1 
assign Y[4'b1011] [59] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^60 ) )   n = 60   d_n = -1 
assign Y[4'b1011] [60] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^61 ) )   n = 61   d_n = -1 
assign Y[4'b1011] [61] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^62 ) )   n = 62   d_n = -1 
assign Y[4'b1011] [62] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^63 ) )   n = 63   d_n = -1 
assign Y[4'b1011] [63] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^64 ) )   n = 64   d_n = -1 
assign Y[4'b1100] [00] = 146'h 000000C041110C4C101000000000000000000;  // -0.4636476090008061 = -1 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = -0-1i 
assign Y[4'b1100] [01] = 146'h 0000003001104101100200000000000000000;  // -0.2449786631268641 = -1 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = -0-1i 
assign Y[4'b1100] [02] = 146'h 0000000C000444104CCC00000000000000000;  // -0.1243549945467614 = -1 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = -0-1i 
assign Y[4'b1100] [03] = 146'h 0000000300001111040420000000000000000;  // -0.0624188099959574 = -1 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = -0-1i 
assign Y[4'b1100] [04] = 146'h 00000000C0000044444100000000000000000;  // -0.0312398334302683 = -1 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = -0-1i 
assign Y[4'b1100] [05] = 146'h 0000000030000001111110000000000000000;  // -0.0156237286204768 = -1 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = -0-1i 
assign Y[4'b1100] [06] = 146'h 000000000C000000044444800000000000000;  // -0.0078123410601011 = -1 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = -0-1i 
assign Y[4'b1100] [07] = 146'h 0000000003000000001111200000000000000;  // -0.0039062301319670 = -1 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = -0-1i 
assign Y[4'b1100] [08] = 146'h 0000000000C00000000044480000000000000;  // -0.0019531225164788 = -1 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = -0-1i 
assign Y[4'b1100] [09] = 146'h 0000000000300000000001120000000000000;  // -0.0009765621895593 = -1 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = -0-1i 
assign Y[4'b1100] [10] = 146'h 00000000000C0000000000048000000000000;  // -0.0004882812111949 = -1 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = -0-1i 
assign Y[4'b1100] [11] = 146'h 0000000000030000000000002000000000000;  // -0.0002441406201494 = -1 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = -0-1i 
assign Y[4'b1100] [12] = 146'h 000000000000C000000000000000000000000;  // -0.0001220703118937 = -1 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = -0-1i 
assign Y[4'b1100] [13] = 146'h 0000000000003000000000000000000000000;  // -0.0000610351561742 = -1 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = -0-1i 
assign Y[4'b1100] [14] = 146'h 0000000000000C00000000000000000000000;  // -0.0000305175781155 = -1 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = -0-1i 
assign Y[4'b1100] [15] = 146'h 0000000000000300000000000000000000000;  // -0.0000152587890613 = -1 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = -0-1i 
assign Y[4'b1100] [16] = 146'h 00000000000000C0000000000000000000000;  // -0.0000076293945311 = -1 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = -0-1i 
assign Y[4'b1100] [17] = 146'h 0000000000000030000000000000000000000;  // -0.0000038146972656 = -1 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = -0-1i 
assign Y[4'b1100] [18] = 146'h 000000000000000C000000000000000000000;  // -0.0000019073486328 = -1 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = -0-1i 
assign Y[4'b1100] [19] = 146'h 0000000000000003000000000000000000000;  // -0.0000009536743164 = -1 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = -0-1i 
assign Y[4'b1100] [20] = 146'h 0000000000000000C00000000000000000000;  // -0.0000004768371582 = -1 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = -0-1i 
assign Y[4'b1100] [21] = 146'h 0000000000000000300000000000000000000;  // -0.0000002384185791 = -1 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = -0-1i 
assign Y[4'b1100] [22] = 146'h 00000000000000000C0000000000000000000;  // -0.0000001192092896 = -1 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = -0-1i 
assign Y[4'b1100] [23] = 146'h 0000000000000000030000000000000000000;  // -0.0000000596046448 = -1 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = -0-1i 
assign Y[4'b1100] [24] = 146'h 000000000000000000C000000000000000000;  // -0.0000000298023224 = -1 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = -0-1i 
assign Y[4'b1100] [25] = 146'h 0000000000000000003000000000000000000;  // -0.0000000149011612 = -1 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = -0-1i 
assign Y[4'b1100] [26] = 146'h 0000000000000000000C00000000000000000;  // -0.0000000074505806 = -1 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = -0-1i 
assign Y[4'b1100] [27] = 146'h 0000000000000000000300000000000000000;  // -0.0000000037252903 = -1 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = -0-1i 
assign Y[4'b1100] [28] = 146'h 00000000000000000000C0000000000000000;  // -0.0000000018626451 = -1 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = -0-1i 
assign Y[4'b1100] [29] = 146'h 0000000000000000000030000000000000000;  // -0.0000000009313226 = -1 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = -0-1i 
assign Y[4'b1100] [30] = 146'h 000000000000000000000C000000000000000;  // -0.0000000004656613 = -1 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = -0-1i 
assign Y[4'b1100] [31] = 146'h 0000000000000000000003000000000000000;  // -0.0000000002328306 = -1 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = -0-1i 
assign Y[4'b1100] [32] = 146'h 0000000000000000000000C00000000000000;  // -0.0000000001164153 = -1 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = -0-1i 
assign Y[4'b1100] [33] = 146'h 0000000000000000000000300000000000000;  // -0.0000000000582077 = -1 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = -0-1i 
assign Y[4'b1100] [34] = 146'h 00000000000000000000000C0000000000000;  // -0.0000000000291038 = -1 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = -0-1i 
assign Y[4'b1100] [35] = 146'h 0000000000000000000000030000000000000;  // -0.0000000000145519 = -1 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = -0-1i 
assign Y[4'b1100] [36] = 146'h 000000000000000000000000C000000000000;  // -0.0000000000072760 = -1 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = -0-1i 
assign Y[4'b1100] [37] = 146'h 0000000000000000000000003000000000000;  // -0.0000000000036380 = -1 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = -0-1i 
assign Y[4'b1100] [38] = 146'h 0000000000000000000000000C00000000000;  // -0.0000000000018190 = -1 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = -0-1i 
assign Y[4'b1100] [39] = 146'h 0000000000000000000000000300000000000;  // -0.0000000000009095 = -1 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = -0-1i 
assign Y[4'b1100] [40] = 146'h 00000000000000000000000000C0000000000;  // -0.0000000000004547 = -1 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = -0-1i 
assign Y[4'b1100] [41] = 146'h 0000000000000000000000000030000000000;  // -0.0000000000002274 = -1 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = -0-1i 
assign Y[4'b1100] [42] = 146'h 000000000000000000000000000C000000000;  // -0.0000000000001137 = -1 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = -0-1i 
assign Y[4'b1100] [43] = 146'h 0000000000000000000000000003000000000;  // -0.0000000000000568 = -1 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = -0-1i 
assign Y[4'b1100] [44] = 146'h 0000000000000000000000000000C00000000;  // -0.0000000000000284 = -1 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = -0-1i 
assign Y[4'b1100] [45] = 146'h 0000000000000000000000000000300000000;  // -0.0000000000000142 = -1 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = -0-1i 
assign Y[4'b1100] [46] = 146'h 00000000000000000000000000000C0000000;  // -0.0000000000000071 = -1 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = -0-1i 
assign Y[4'b1100] [47] = 146'h 0000000000000000000000000000030000000;  // -0.0000000000000036 = -1 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = -0-1i 
assign Y[4'b1100] [48] = 146'h 000000000000000000000000000000C000000;  // -0.0000000000000018 = -1 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = -0-1i 
assign Y[4'b1100] [49] = 146'h 0000000000000000000000000000003000000;  // -0.0000000000000009 = -1 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = -0-1i 
assign Y[4'b1100] [50] = 146'h 0000000000000000000000000000000C00000;  // -0.0000000000000004 = -1 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = -0-1i 
assign Y[4'b1100] [51] = 146'h 0000000000000000000000000000000300000;  // -0.0000000000000002 = -1 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = -0-1i 
assign Y[4'b1100] [52] = 146'h 00000000000000000000000000000000C0000;  // -0.0000000000000001 = -1 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = -0-1i 
assign Y[4'b1100] [53] = 146'h 0000000000000000000000000000000030000;  // -0.0000000000000001 = -1 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = -0-1i 
assign Y[4'b1100] [54] = 146'h 000000000000000000000000000000000C000;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = -0-1i 
assign Y[4'b1100] [55] = 146'h 0000000000000000000000000000000003000;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = -0-1i 
assign Y[4'b1100] [56] = 146'h 0000000000000000000000000000000000C00;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = -0-1i 
assign Y[4'b1100] [57] = 146'h 0000000000000000000000000000000000300;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = -0-1i 
assign Y[4'b1100] [58] = 146'h 00000000000000000000000000000000000C0;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = -0-1i 
assign Y[4'b1100] [59] = 146'h 0000000000000000000000000000000000030;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = -0-1i 
assign Y[4'b1100] [60] = 146'h 000000000000000000000000000000000000C;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = -0-1i 
assign Y[4'b1100] [61] = 146'h 0000000000000000000000000000000000003;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = -0-1i 
assign Y[4'b1100] [62] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = -0-1i 
assign Y[4'b1100] [63] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = -0-1i 
assign Y[4'b1101] [00] = 146'h 000000330CC4043004C400000000000000000;  // -0.3217505543966422 = -1 * atan( 1 / (  1 + 2^1 ) )   n =  1   d_n = 1-1i 
assign Y[4'b1101] [01] = 146'h 000000310CC0C0C0300200000000000000000;  // -0.1973955598498807 = -1 * atan( 1 / (  1 + 2^2 ) )   n =  2   d_n = 1-1i 
assign Y[4'b1101] [02] = 146'h 0000000C10333000C00C80000000000000000;  // -0.1106572211738956 = -1 * atan( 1 / (  1 + 2^3 ) )   n =  3   d_n = 1-1i 
assign Y[4'b1101] [03] = 146'h 000000030100CCCC010C00000000000000000;  // -0.0587558227157227 = -1 * atan( 1 / (  1 + 2^4 ) )   n =  4   d_n = 1-1i 
assign Y[4'b1101] [04] = 146'h 00000000C0100333330130000000000000000;  // -0.0302937599187751 = -1 * atan( 1 / (  1 + 2^5 ) )   n =  5   d_n = 1-1i 
assign Y[4'b1101] [05] = 146'h 000000003001000CCCCCC0000000000000000;  // -0.0153834017805952 = -1 * atan( 1 / (  1 + 2^6 ) )   n =  6   d_n = 1-1i 
assign Y[4'b1101] [06] = 146'h 000000000C001000333333000000000000000;  // -0.0077517827122069 = -1 * atan( 1 / (  1 + 2^7 ) )   n =  7   d_n = 1-1i 
assign Y[4'b1101] [07] = 146'h 000000000300010000CCCCC00000000000000;  // -0.0038910309466445 = -1 * atan( 1 / (  1 + 2^8 ) )   n =  8   d_n = 1-1i 
assign Y[4'b1101] [08] = 146'h 0000000000C00010000333300000000000000;  // -0.0019493152697654 = -1 * atan( 1 / (  1 + 2^9 ) )   n =  9   d_n = 1-1i 
assign Y[4'b1101] [09] = 146'h 000000000030000100000CCC0000000000000;  // -0.0009756094465646 = -1 * atan( 1 / (  1 + 2^10 ) )   n = 10   d_n = 1-1i 
assign Y[4'b1101] [10] = 146'h 00000000000C0000100000330000000000000;  // -0.0004880429090311 = -1 * atan( 1 / (  1 + 2^11 ) )   n = 11   d_n = 1-1i 
assign Y[4'b1101] [11] = 146'h 000000000003000001000000C000000000000;  // -0.0002440810300565 = -1 * atan( 1 / (  1 + 2^12 ) )   n = 12   d_n = 1-1i 
assign Y[4'b1101] [12] = 146'h 000000000000C000001000000000000000000;  // -0.0001220554125515 = -1 * atan( 1 / (  1 + 2^13 ) )   n = 13   d_n = 1-1i 
assign Y[4'b1101] [13] = 146'h 0000000000003000000100000000000000000;  // -0.0000610314311113 = -1 * atan( 1 / (  1 + 2^14 ) )   n = 14   d_n = 1-1i 
assign Y[4'b1101] [14] = 146'h 0000000000000C00000010000000000000000;  // -0.0000305166468214 = -1 * atan( 1 / (  1 + 2^15 ) )   n = 15   d_n = 1-1i 
assign Y[4'b1101] [15] = 146'h 0000000000000300000001000000000000000;  // -0.0000152585562342 = -1 * atan( 1 / (  1 + 2^16 ) )   n = 16   d_n = 1-1i 
assign Y[4'b1101] [16] = 146'h 00000000000000C0000000100000000000000;  // -0.0000076293363239 = -1 * atan( 1 / (  1 + 2^17 ) )   n = 17   d_n = 1-1i 
assign Y[4'b1101] [17] = 146'h 0000000000000030000000010000000000000;  // -0.0000038146827137 = -1 * atan( 1 / (  1 + 2^18 ) )   n = 18   d_n = 1-1i 
assign Y[4'b1101] [18] = 146'h 000000000000000C000000001000000000000;  // -0.0000019073449948 = -1 * atan( 1 / (  1 + 2^19 ) )   n = 19   d_n = 1-1i 
assign Y[4'b1101] [19] = 146'h 0000000000000003000000000100000000000;  // -0.0000009536734069 = -1 * atan( 1 / (  1 + 2^20 ) )   n = 20   d_n = 1-1i 
assign Y[4'b1101] [20] = 146'h 0000000000000000C00000000010000000000;  // -0.0000004768369308 = -1 * atan( 1 / (  1 + 2^21 ) )   n = 21   d_n = 1-1i 
assign Y[4'b1101] [21] = 146'h 0000000000000000300000000001000000000;  // -0.0000002384185223 = -1 * atan( 1 / (  1 + 2^22 ) )   n = 22   d_n = 1-1i 
assign Y[4'b1101] [22] = 146'h 00000000000000000C0000000000100000000;  // -0.0000001192092753 = -1 * atan( 1 / (  1 + 2^23 ) )   n = 23   d_n = 1-1i 
assign Y[4'b1101] [23] = 146'h 0000000000000000030000000000010000000;  // -0.0000000596046412 = -1 * atan( 1 / (  1 + 2^24 ) )   n = 24   d_n = 1-1i 
assign Y[4'b1101] [24] = 146'h 000000000000000000C000000000001000000;  // -0.0000000298023215 = -1 * atan( 1 / (  1 + 2^25 ) )   n = 25   d_n = 1-1i 
assign Y[4'b1101] [25] = 146'h 0000000000000000003000000000000000000;  // -0.0000000149011610 = -1 * atan( 1 / (  1 + 2^26 ) )   n = 26   d_n = 1-1i 
assign Y[4'b1101] [26] = 146'h 0000000000000000000C00000000000000000;  // -0.0000000074505805 = -1 * atan( 1 / (  1 + 2^27 ) )   n = 27   d_n = 1-1i 
assign Y[4'b1101] [27] = 146'h 0000000000000000000300000000000000000;  // -0.0000000037252903 = -1 * atan( 1 / (  1 + 2^28 ) )   n = 28   d_n = 1-1i 
assign Y[4'b1101] [28] = 146'h 00000000000000000000C0000000000000000;  // -0.0000000018626451 = -1 * atan( 1 / (  1 + 2^29 ) )   n = 29   d_n = 1-1i 
assign Y[4'b1101] [29] = 146'h 0000000000000000000030000000000000000;  // -0.0000000009313226 = -1 * atan( 1 / (  1 + 2^30 ) )   n = 30   d_n = 1-1i 
assign Y[4'b1101] [30] = 146'h 000000000000000000000C000000000000000;  // -0.0000000004656613 = -1 * atan( 1 / (  1 + 2^31 ) )   n = 31   d_n = 1-1i 
assign Y[4'b1101] [31] = 146'h 0000000000000000000003000000000000000;  // -0.0000000002328306 = -1 * atan( 1 / (  1 + 2^32 ) )   n = 32   d_n = 1-1i 
assign Y[4'b1101] [32] = 146'h 0000000000000000000000C00000000000000;  // -0.0000000001164153 = -1 * atan( 1 / (  1 + 2^33 ) )   n = 33   d_n = 1-1i 
assign Y[4'b1101] [33] = 146'h 0000000000000000000000300000000000000;  // -0.0000000000582077 = -1 * atan( 1 / (  1 + 2^34 ) )   n = 34   d_n = 1-1i 
assign Y[4'b1101] [34] = 146'h 00000000000000000000000C0000000000000;  // -0.0000000000291038 = -1 * atan( 1 / (  1 + 2^35 ) )   n = 35   d_n = 1-1i 
assign Y[4'b1101] [35] = 146'h 0000000000000000000000030000000000000;  // -0.0000000000145519 = -1 * atan( 1 / (  1 + 2^36 ) )   n = 36   d_n = 1-1i 
assign Y[4'b1101] [36] = 146'h 000000000000000000000000C000000000000;  // -0.0000000000072760 = -1 * atan( 1 / (  1 + 2^37 ) )   n = 37   d_n = 1-1i 
assign Y[4'b1101] [37] = 146'h 0000000000000000000000003000000000000;  // -0.0000000000036380 = -1 * atan( 1 / (  1 + 2^38 ) )   n = 38   d_n = 1-1i 
assign Y[4'b1101] [38] = 146'h 0000000000000000000000000C00000000000;  // -0.0000000000018190 = -1 * atan( 1 / (  1 + 2^39 ) )   n = 39   d_n = 1-1i 
assign Y[4'b1101] [39] = 146'h 0000000000000000000000000300000000000;  // -0.0000000000009095 = -1 * atan( 1 / (  1 + 2^40 ) )   n = 40   d_n = 1-1i 
assign Y[4'b1101] [40] = 146'h 00000000000000000000000000C0000000000;  // -0.0000000000004547 = -1 * atan( 1 / (  1 + 2^41 ) )   n = 41   d_n = 1-1i 
assign Y[4'b1101] [41] = 146'h 0000000000000000000000000030000000000;  // -0.0000000000002274 = -1 * atan( 1 / (  1 + 2^42 ) )   n = 42   d_n = 1-1i 
assign Y[4'b1101] [42] = 146'h 000000000000000000000000000C000000000;  // -0.0000000000001137 = -1 * atan( 1 / (  1 + 2^43 ) )   n = 43   d_n = 1-1i 
assign Y[4'b1101] [43] = 146'h 0000000000000000000000000003000000000;  // -0.0000000000000568 = -1 * atan( 1 / (  1 + 2^44 ) )   n = 44   d_n = 1-1i 
assign Y[4'b1101] [44] = 146'h 0000000000000000000000000000C00000000;  // -0.0000000000000284 = -1 * atan( 1 / (  1 + 2^45 ) )   n = 45   d_n = 1-1i 
assign Y[4'b1101] [45] = 146'h 0000000000000000000000000000300000000;  // -0.0000000000000142 = -1 * atan( 1 / (  1 + 2^46 ) )   n = 46   d_n = 1-1i 
assign Y[4'b1101] [46] = 146'h 00000000000000000000000000000C0000000;  // -0.0000000000000071 = -1 * atan( 1 / (  1 + 2^47 ) )   n = 47   d_n = 1-1i 
assign Y[4'b1101] [47] = 146'h 0000000000000000000000000000030000000;  // -0.0000000000000036 = -1 * atan( 1 / (  1 + 2^48 ) )   n = 48   d_n = 1-1i 
assign Y[4'b1101] [48] = 146'h 000000000000000000000000000000C000000;  // -0.0000000000000018 = -1 * atan( 1 / (  1 + 2^49 ) )   n = 49   d_n = 1-1i 
assign Y[4'b1101] [49] = 146'h 0000000000000000000000000000003000000;  // -0.0000000000000009 = -1 * atan( 1 / (  1 + 2^50 ) )   n = 50   d_n = 1-1i 
assign Y[4'b1101] [50] = 146'h 0000000000000000000000000000000C00000;  // -0.0000000000000004 = -1 * atan( 1 / (  1 + 2^51 ) )   n = 51   d_n = 1-1i 
assign Y[4'b1101] [51] = 146'h 0000000000000000000000000000000300000;  // -0.0000000000000002 = -1 * atan( 1 / (  1 + 2^52 ) )   n = 52   d_n = 1-1i 
assign Y[4'b1101] [52] = 146'h 00000000000000000000000000000000C0000;  // -0.0000000000000001 = -1 * atan( 1 / (  1 + 2^53 ) )   n = 53   d_n = 1-1i 
assign Y[4'b1101] [53] = 146'h 0000000000000000000000000000000030000;  // -0.0000000000000001 = -1 * atan( 1 / (  1 + 2^54 ) )   n = 54   d_n = 1-1i 
assign Y[4'b1101] [54] = 146'h 000000000000000000000000000000000C000;  // -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^55 ) )   n = 55   d_n = 1-1i 
assign Y[4'b1101] [55] = 146'h 0000000000000000000000000000000003000;  // -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^56 ) )   n = 56   d_n = 1-1i 
assign Y[4'b1101] [56] = 146'h 0000000000000000000000000000000000C00;  // -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^57 ) )   n = 57   d_n = 1-1i 
assign Y[4'b1101] [57] = 146'h 0000000000000000000000000000000000300;  // -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^58 ) )   n = 58   d_n = 1-1i 
assign Y[4'b1101] [58] = 146'h 00000000000000000000000000000000000C0;  // -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^59 ) )   n = 59   d_n = 1-1i 
assign Y[4'b1101] [59] = 146'h 0000000000000000000000000000000000030;  // -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^60 ) )   n = 60   d_n = 1-1i 
assign Y[4'b1101] [60] = 146'h 000000000000000000000000000000000000C;  // -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^61 ) )   n = 61   d_n = 1-1i 
assign Y[4'b1101] [61] = 146'h 0000000000000000000000000000000000003;  // -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^62 ) )   n = 62   d_n = 1-1i 
assign Y[4'b1101] [62] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^63 ) )   n = 63   d_n = 1-1i 
assign Y[4'b1101] [63] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^64 ) )   n = 64   d_n = 1-1i 
assign Y[4'b1110] [00] = 146'h 000000C041110C4C101000000000000000000;  // -0.4636476090008061 = -1 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = -0-1i 
assign Y[4'b1110] [01] = 146'h 0000003001104101100200000000000000000;  // -0.2449786631268641 = -1 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = -0-1i 
assign Y[4'b1110] [02] = 146'h 0000000C000444104CCC00000000000000000;  // -0.1243549945467614 = -1 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = -0-1i 
assign Y[4'b1110] [03] = 146'h 0000000300001111040420000000000000000;  // -0.0624188099959574 = -1 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = -0-1i 
assign Y[4'b1110] [04] = 146'h 00000000C0000044444100000000000000000;  // -0.0312398334302683 = -1 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = -0-1i 
assign Y[4'b1110] [05] = 146'h 0000000030000001111110000000000000000;  // -0.0156237286204768 = -1 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = -0-1i 
assign Y[4'b1110] [06] = 146'h 000000000C000000044444800000000000000;  // -0.0078123410601011 = -1 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = -0-1i 
assign Y[4'b1110] [07] = 146'h 0000000003000000001111200000000000000;  // -0.0039062301319670 = -1 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = -0-1i 
assign Y[4'b1110] [08] = 146'h 0000000000C00000000044480000000000000;  // -0.0019531225164788 = -1 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = -0-1i 
assign Y[4'b1110] [09] = 146'h 0000000000300000000001120000000000000;  // -0.0009765621895593 = -1 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = -0-1i 
assign Y[4'b1110] [10] = 146'h 00000000000C0000000000048000000000000;  // -0.0004882812111949 = -1 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = -0-1i 
assign Y[4'b1110] [11] = 146'h 0000000000030000000000002000000000000;  // -0.0002441406201494 = -1 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = -0-1i 
assign Y[4'b1110] [12] = 146'h 000000000000C000000000000000000000000;  // -0.0001220703118937 = -1 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = -0-1i 
assign Y[4'b1110] [13] = 146'h 0000000000003000000000000000000000000;  // -0.0000610351561742 = -1 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = -0-1i 
assign Y[4'b1110] [14] = 146'h 0000000000000C00000000000000000000000;  // -0.0000305175781155 = -1 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = -0-1i 
assign Y[4'b1110] [15] = 146'h 0000000000000300000000000000000000000;  // -0.0000152587890613 = -1 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = -0-1i 
assign Y[4'b1110] [16] = 146'h 00000000000000C0000000000000000000000;  // -0.0000076293945311 = -1 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = -0-1i 
assign Y[4'b1110] [17] = 146'h 0000000000000030000000000000000000000;  // -0.0000038146972656 = -1 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = -0-1i 
assign Y[4'b1110] [18] = 146'h 000000000000000C000000000000000000000;  // -0.0000019073486328 = -1 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = -0-1i 
assign Y[4'b1110] [19] = 146'h 0000000000000003000000000000000000000;  // -0.0000009536743164 = -1 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = -0-1i 
assign Y[4'b1110] [20] = 146'h 0000000000000000C00000000000000000000;  // -0.0000004768371582 = -1 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = -0-1i 
assign Y[4'b1110] [21] = 146'h 0000000000000000300000000000000000000;  // -0.0000002384185791 = -1 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = -0-1i 
assign Y[4'b1110] [22] = 146'h 00000000000000000C0000000000000000000;  // -0.0000001192092896 = -1 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = -0-1i 
assign Y[4'b1110] [23] = 146'h 0000000000000000030000000000000000000;  // -0.0000000596046448 = -1 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = -0-1i 
assign Y[4'b1110] [24] = 146'h 000000000000000000C000000000000000000;  // -0.0000000298023224 = -1 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = -0-1i 
assign Y[4'b1110] [25] = 146'h 0000000000000000003000000000000000000;  // -0.0000000149011612 = -1 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = -0-1i 
assign Y[4'b1110] [26] = 146'h 0000000000000000000C00000000000000000;  // -0.0000000074505806 = -1 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = -0-1i 
assign Y[4'b1110] [27] = 146'h 0000000000000000000300000000000000000;  // -0.0000000037252903 = -1 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = -0-1i 
assign Y[4'b1110] [28] = 146'h 00000000000000000000C0000000000000000;  // -0.0000000018626451 = -1 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = -0-1i 
assign Y[4'b1110] [29] = 146'h 0000000000000000000030000000000000000;  // -0.0000000009313226 = -1 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = -0-1i 
assign Y[4'b1110] [30] = 146'h 000000000000000000000C000000000000000;  // -0.0000000004656613 = -1 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = -0-1i 
assign Y[4'b1110] [31] = 146'h 0000000000000000000003000000000000000;  // -0.0000000002328306 = -1 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = -0-1i 
assign Y[4'b1110] [32] = 146'h 0000000000000000000000C00000000000000;  // -0.0000000001164153 = -1 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = -0-1i 
assign Y[4'b1110] [33] = 146'h 0000000000000000000000300000000000000;  // -0.0000000000582077 = -1 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = -0-1i 
assign Y[4'b1110] [34] = 146'h 00000000000000000000000C0000000000000;  // -0.0000000000291038 = -1 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = -0-1i 
assign Y[4'b1110] [35] = 146'h 0000000000000000000000030000000000000;  // -0.0000000000145519 = -1 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = -0-1i 
assign Y[4'b1110] [36] = 146'h 000000000000000000000000C000000000000;  // -0.0000000000072760 = -1 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = -0-1i 
assign Y[4'b1110] [37] = 146'h 0000000000000000000000003000000000000;  // -0.0000000000036380 = -1 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = -0-1i 
assign Y[4'b1110] [38] = 146'h 0000000000000000000000000C00000000000;  // -0.0000000000018190 = -1 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = -0-1i 
assign Y[4'b1110] [39] = 146'h 0000000000000000000000000300000000000;  // -0.0000000000009095 = -1 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = -0-1i 
assign Y[4'b1110] [40] = 146'h 00000000000000000000000000C0000000000;  // -0.0000000000004547 = -1 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = -0-1i 
assign Y[4'b1110] [41] = 146'h 0000000000000000000000000030000000000;  // -0.0000000000002274 = -1 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = -0-1i 
assign Y[4'b1110] [42] = 146'h 000000000000000000000000000C000000000;  // -0.0000000000001137 = -1 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = -0-1i 
assign Y[4'b1110] [43] = 146'h 0000000000000000000000000003000000000;  // -0.0000000000000568 = -1 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = -0-1i 
assign Y[4'b1110] [44] = 146'h 0000000000000000000000000000C00000000;  // -0.0000000000000284 = -1 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = -0-1i 
assign Y[4'b1110] [45] = 146'h 0000000000000000000000000000300000000;  // -0.0000000000000142 = -1 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = -0-1i 
assign Y[4'b1110] [46] = 146'h 00000000000000000000000000000C0000000;  // -0.0000000000000071 = -1 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = -0-1i 
assign Y[4'b1110] [47] = 146'h 0000000000000000000000000000030000000;  // -0.0000000000000036 = -1 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = -0-1i 
assign Y[4'b1110] [48] = 146'h 000000000000000000000000000000C000000;  // -0.0000000000000018 = -1 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = -0-1i 
assign Y[4'b1110] [49] = 146'h 0000000000000000000000000000003000000;  // -0.0000000000000009 = -1 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = -0-1i 
assign Y[4'b1110] [50] = 146'h 0000000000000000000000000000000C00000;  // -0.0000000000000004 = -1 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = -0-1i 
assign Y[4'b1110] [51] = 146'h 0000000000000000000000000000000300000;  // -0.0000000000000002 = -1 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = -0-1i 
assign Y[4'b1110] [52] = 146'h 00000000000000000000000000000000C0000;  // -0.0000000000000001 = -1 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = -0-1i 
assign Y[4'b1110] [53] = 146'h 0000000000000000000000000000000030000;  // -0.0000000000000001 = -1 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = -0-1i 
assign Y[4'b1110] [54] = 146'h 000000000000000000000000000000000C000;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = -0-1i 
assign Y[4'b1110] [55] = 146'h 0000000000000000000000000000000003000;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = -0-1i 
assign Y[4'b1110] [56] = 146'h 0000000000000000000000000000000000C00;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = -0-1i 
assign Y[4'b1110] [57] = 146'h 0000000000000000000000000000000000300;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = -0-1i 
assign Y[4'b1110] [58] = 146'h 00000000000000000000000000000000000C0;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = -0-1i 
assign Y[4'b1110] [59] = 146'h 0000000000000000000000000000000000030;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = -0-1i 
assign Y[4'b1110] [60] = 146'h 000000000000000000000000000000000000C;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = -0-1i 
assign Y[4'b1110] [61] = 146'h 0000000000000000000000000000000000003;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = -0-1i 
assign Y[4'b1110] [62] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = -0-1i 
assign Y[4'b1110] [63] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = -0-1i 
assign Y[4'b1111] [00] = 146'h 00000310C30300044CC000000000000000000;  // -0.7853981633974483 = -1 * atan( 1 / ( -1 + 2^1 ) )   n =  1   d_n = -1-1i 
assign Y[4'b1111] [01] = 146'h 000000330CC4043004C400000000000000000;  // -0.3217505543966422 = -1 * atan( 1 / ( -1 + 2^2 ) )   n =  2   d_n = -1-1i 
assign Y[4'b1111] [02] = 146'h 0000000C30333044044100000000000000000;  // -0.1418970546041639 = -1 * atan( 1 / ( -1 + 2^3 ) )   n =  3   d_n = -1-1i 
assign Y[4'b1111] [03] = 146'h 000000030300CCCC10C040000000000000000;  // -0.0665681637758238 = -1 * atan( 1 / ( -1 + 2^4 ) )   n =  4   d_n = -1-1i 
assign Y[4'b1111] [04] = 146'h 00000000C03003333304D0000000000000000;  // -0.0322468824352539 = -1 * atan( 1 / ( -1 + 2^5 ) )   n =  5   d_n = -1-1i 
assign Y[4'b1111] [05] = 146'h 000000003003000CCCCCC0000000000000000;  // -0.0158716829917901 = -1 * atan( 1 / ( -1 + 2^6 ) )   n =  6   d_n = -1-1i 
assign Y[4'b1111] [06] = 146'h 000000000C003000333333000000000000000;  // -0.0078738530241005 = -1 * atan( 1 / ( -1 + 2^7 ) )   n =  7   d_n = -1-1i 
assign Y[4'b1111] [07] = 146'h 000000000300030000CCCCC00000000000000;  // -0.0039215485247600 = -1 * atan( 1 / ( -1 + 2^8 ) )   n =  8   d_n = -1-1i 
assign Y[4'b1111] [08] = 146'h 0000000000C00030000333300000000000000;  // -0.0019569446642965 = -1 * atan( 1 / ( -1 + 2^9 ) )   n =  9   d_n = -1-1i 
assign Y[4'b1111] [09] = 146'h 000000000030000300000CCC0000000000000;  // -0.0009775167951974 = -1 * atan( 1 / ( -1 + 2^10 ) )   n = 10   d_n = -1-1i 
assign Y[4'b1111] [10] = 146'h 00000000000C0000300000330000000000000;  // -0.0004885197461893 = -1 * atan( 1 / ( -1 + 2^11 ) )   n = 11   d_n = -1-1i 
assign Y[4'b1111] [11] = 146'h 000000000003000003000000C000000000000;  // -0.0002442002393461 = -1 * atan( 1 / ( -1 + 2^12 ) )   n = 12   d_n = -1-1i 
assign Y[4'b1111] [12] = 146'h 000000000000C000003000000000000000000;  // -0.0001220852148739 = -1 * atan( 1 / ( -1 + 2^13 ) )   n = 13   d_n = -1-1i 
assign Y[4'b1111] [13] = 146'h 0000000000003000000300000000000000000;  // -0.0000610388816919 = -1 * atan( 1 / ( -1 + 2^14 ) )   n = 14   d_n = -1-1i 
assign Y[4'b1111] [14] = 146'h 0000000000000C00000030000000000000000;  // -0.0000305185094665 = -1 * atan( 1 / ( -1 + 2^15 ) )   n = 15   d_n = -1-1i 
assign Y[4'b1111] [15] = 146'h 0000000000000300000003000000000000000;  // -0.0000152590218955 = -1 * atan( 1 / ( -1 + 2^16 ) )   n = 16   d_n = -1-1i 
assign Y[4'b1111] [16] = 146'h 00000000000000C0000000300000000000000;  // -0.0000076294527392 = -1 * atan( 1 / ( -1 + 2^17 ) )   n = 17   d_n = -1-1i 
assign Y[4'b1111] [17] = 146'h 0000000000000030000000030000000000000;  // -0.0000038147118176 = -1 * atan( 1 / ( -1 + 2^18 ) )   n = 18   d_n = -1-1i 
assign Y[4'b1111] [18] = 146'h 000000000000000C000000003000000000000;  // -0.0000019073522708 = -1 * atan( 1 / ( -1 + 2^19 ) )   n = 19   d_n = -1-1i 
assign Y[4'b1111] [19] = 146'h 0000000000000003000000000300000000000;  // -0.0000009536752259 = -1 * atan( 1 / ( -1 + 2^20 ) )   n = 20   d_n = -1-1i 
assign Y[4'b1111] [20] = 146'h 0000000000000000C00000000030000000000;  // -0.0000004768373856 = -1 * atan( 1 / ( -1 + 2^21 ) )   n = 21   d_n = -1-1i 
assign Y[4'b1111] [21] = 146'h 0000000000000000300000000003000000000;  // -0.0000002384186359 = -1 * atan( 1 / ( -1 + 2^22 ) )   n = 22   d_n = -1-1i 
assign Y[4'b1111] [22] = 146'h 00000000000000000C0000000000300000000;  // -0.0000001192093038 = -1 * atan( 1 / ( -1 + 2^23 ) )   n = 23   d_n = -1-1i 
assign Y[4'b1111] [23] = 146'h 0000000000000000030000000000030000000;  // -0.0000000596046483 = -1 * atan( 1 / ( -1 + 2^24 ) )   n = 24   d_n = -1-1i 
assign Y[4'b1111] [24] = 146'h 000000000000000000C000000000003000000;  // -0.0000000298023233 = -1 * atan( 1 / ( -1 + 2^25 ) )   n = 25   d_n = -1-1i 
assign Y[4'b1111] [25] = 146'h 0000000000000000003000000000000400000;  // -0.0000000149011614 = -1 * atan( 1 / ( -1 + 2^26 ) )   n = 26   d_n = -1-1i 
assign Y[4'b1111] [26] = 146'h 0000000000000000000C00000000000000000;  // -0.0000000074505807 = -1 * atan( 1 / ( -1 + 2^27 ) )   n = 27   d_n = -1-1i 
assign Y[4'b1111] [27] = 146'h 0000000000000000000300000000000000000;  // -0.0000000037252903 = -1 * atan( 1 / ( -1 + 2^28 ) )   n = 28   d_n = -1-1i 
assign Y[4'b1111] [28] = 146'h 00000000000000000000C0000000000000000;  // -0.0000000018626452 = -1 * atan( 1 / ( -1 + 2^29 ) )   n = 29   d_n = -1-1i 
assign Y[4'b1111] [29] = 146'h 0000000000000000000030000000000000000;  // -0.0000000009313226 = -1 * atan( 1 / ( -1 + 2^30 ) )   n = 30   d_n = -1-1i 
assign Y[4'b1111] [30] = 146'h 000000000000000000000C000000000000000;  // -0.0000000004656613 = -1 * atan( 1 / ( -1 + 2^31 ) )   n = 31   d_n = -1-1i 
assign Y[4'b1111] [31] = 146'h 0000000000000000000003000000000000000;  // -0.0000000002328306 = -1 * atan( 1 / ( -1 + 2^32 ) )   n = 32   d_n = -1-1i 
assign Y[4'b1111] [32] = 146'h 0000000000000000000000C00000000000000;  // -0.0000000001164153 = -1 * atan( 1 / ( -1 + 2^33 ) )   n = 33   d_n = -1-1i 
assign Y[4'b1111] [33] = 146'h 0000000000000000000000300000000000000;  // -0.0000000000582077 = -1 * atan( 1 / ( -1 + 2^34 ) )   n = 34   d_n = -1-1i 
assign Y[4'b1111] [34] = 146'h 00000000000000000000000C0000000000000;  // -0.0000000000291038 = -1 * atan( 1 / ( -1 + 2^35 ) )   n = 35   d_n = -1-1i 
assign Y[4'b1111] [35] = 146'h 0000000000000000000000030000000000000;  // -0.0000000000145519 = -1 * atan( 1 / ( -1 + 2^36 ) )   n = 36   d_n = -1-1i 
assign Y[4'b1111] [36] = 146'h 000000000000000000000000C000000000000;  // -0.0000000000072760 = -1 * atan( 1 / ( -1 + 2^37 ) )   n = 37   d_n = -1-1i 
assign Y[4'b1111] [37] = 146'h 0000000000000000000000003000000000000;  // -0.0000000000036380 = -1 * atan( 1 / ( -1 + 2^38 ) )   n = 38   d_n = -1-1i 
assign Y[4'b1111] [38] = 146'h 0000000000000000000000000C00000000000;  // -0.0000000000018190 = -1 * atan( 1 / ( -1 + 2^39 ) )   n = 39   d_n = -1-1i 
assign Y[4'b1111] [39] = 146'h 0000000000000000000000000300000000000;  // -0.0000000000009095 = -1 * atan( 1 / ( -1 + 2^40 ) )   n = 40   d_n = -1-1i 
assign Y[4'b1111] [40] = 146'h 00000000000000000000000000C0000000000;  // -0.0000000000004547 = -1 * atan( 1 / ( -1 + 2^41 ) )   n = 41   d_n = -1-1i 
assign Y[4'b1111] [41] = 146'h 0000000000000000000000000030000000000;  // -0.0000000000002274 = -1 * atan( 1 / ( -1 + 2^42 ) )   n = 42   d_n = -1-1i 
assign Y[4'b1111] [42] = 146'h 000000000000000000000000000C000000000;  // -0.0000000000001137 = -1 * atan( 1 / ( -1 + 2^43 ) )   n = 43   d_n = -1-1i 
assign Y[4'b1111] [43] = 146'h 0000000000000000000000000003000000000;  // -0.0000000000000568 = -1 * atan( 1 / ( -1 + 2^44 ) )   n = 44   d_n = -1-1i 
assign Y[4'b1111] [44] = 146'h 0000000000000000000000000000C00000000;  // -0.0000000000000284 = -1 * atan( 1 / ( -1 + 2^45 ) )   n = 45   d_n = -1-1i 
assign Y[4'b1111] [45] = 146'h 0000000000000000000000000000300000000;  // -0.0000000000000142 = -1 * atan( 1 / ( -1 + 2^46 ) )   n = 46   d_n = -1-1i 
assign Y[4'b1111] [46] = 146'h 00000000000000000000000000000C0000000;  // -0.0000000000000071 = -1 * atan( 1 / ( -1 + 2^47 ) )   n = 47   d_n = -1-1i 
assign Y[4'b1111] [47] = 146'h 0000000000000000000000000000030000000;  // -0.0000000000000036 = -1 * atan( 1 / ( -1 + 2^48 ) )   n = 48   d_n = -1-1i 
assign Y[4'b1111] [48] = 146'h 000000000000000000000000000000C000000;  // -0.0000000000000018 = -1 * atan( 1 / ( -1 + 2^49 ) )   n = 49   d_n = -1-1i 
assign Y[4'b1111] [49] = 146'h 0000000000000000000000000000003000000;  // -0.0000000000000009 = -1 * atan( 1 / ( -1 + 2^50 ) )   n = 50   d_n = -1-1i 
assign Y[4'b1111] [50] = 146'h 0000000000000000000000000000000C00000;  // -0.0000000000000004 = -1 * atan( 1 / ( -1 + 2^51 ) )   n = 51   d_n = -1-1i 
assign Y[4'b1111] [51] = 146'h 0000000000000000000000000000000300000;  // -0.0000000000000002 = -1 * atan( 1 / ( -1 + 2^52 ) )   n = 52   d_n = -1-1i 
assign Y[4'b1111] [52] = 146'h 00000000000000000000000000000000C0000;  // -0.0000000000000001 = -1 * atan( 1 / ( -1 + 2^53 ) )   n = 53   d_n = -1-1i 
assign Y[4'b1111] [53] = 146'h 0000000000000000000000000000000030000;  // -0.0000000000000001 = -1 * atan( 1 / ( -1 + 2^54 ) )   n = 54   d_n = -1-1i 
assign Y[4'b1111] [54] = 146'h 000000000000000000000000000000000C000;  // -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^55 ) )   n = 55   d_n = -1-1i 
assign Y[4'b1111] [55] = 146'h 0000000000000000000000000000000003000;  // -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^56 ) )   n = 56   d_n = -1-1i 
assign Y[4'b1111] [56] = 146'h 0000000000000000000000000000000000C00;  // -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^57 ) )   n = 57   d_n = -1-1i 
assign Y[4'b1111] [57] = 146'h 0000000000000000000000000000000000300;  // -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^58 ) )   n = 58   d_n = -1-1i 
assign Y[4'b1111] [58] = 146'h 00000000000000000000000000000000000C0;  // -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^59 ) )   n = 59   d_n = -1-1i 
assign Y[4'b1111] [59] = 146'h 0000000000000000000000000000000000030;  // -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^60 ) )   n = 60   d_n = -1-1i 
assign Y[4'b1111] [60] = 146'h 000000000000000000000000000000000000C;  // -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^61 ) )   n = 61   d_n = -1-1i 
assign Y[4'b1111] [61] = 146'h 0000000000000000000000000000000000003;  // -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^62 ) )   n = 62   d_n = -1-1i 
assign Y[4'b1111] [62] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^63 ) )   n = 63   d_n = -1-1i 
assign Y[4'b1111] [63] = 146'h 0000000000000000000000000000000000000;  // -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^64 ) )   n = 64   d_n = -1-1i 
assign u[4'b0000] [00] = 21'h 000000;  // +0.0000000000000000 = 2^ 1 * ln( 1 +  0 * 2^(- 1+1) + ( 0^2+ 0^2) * 2^(-2* 1) )   n =  1   d_n = 0 
assign u[4'b0000] [01] = 21'h 000000;  // +0.0000000000000000 = 2^ 2 * ln( 1 +  0 * 2^(- 2+1) + ( 0^2+ 0^2) * 2^(-2* 2) )   n =  2   d_n = 0 
assign u[4'b0000] [02] = 21'h 000000;  // +0.0000000000000000 = 2^ 3 * ln( 1 +  0 * 2^(- 3+1) + ( 0^2+ 0^2) * 2^(-2* 3) )   n =  3   d_n = 0 
assign u[4'b0000] [03] = 21'h 000000;  // +0.0000000000000000 = 2^ 4 * ln( 1 +  0 * 2^(- 4+1) + ( 0^2+ 0^2) * 2^(-2* 4) )   n =  4   d_n = 0 
assign u[4'b0000] [04] = 21'h 000000;  // +0.0000000000000000 = 2^ 5 * ln( 1 +  0 * 2^(- 5+1) + ( 0^2+ 0^2) * 2^(-2* 5) )   n =  5   d_n = 0 
assign u[4'b0000] [05] = 21'h 000000;  // +0.0000000000000000 = 2^ 6 * ln( 1 +  0 * 2^(- 6+1) + ( 0^2+ 0^2) * 2^(-2* 6) )   n =  6   d_n = 0 
assign u[4'b0000] [06] = 21'h 000000;  // +0.0000000000000000 = 2^ 7 * ln( 1 +  0 * 2^(- 7+1) + ( 0^2+ 0^2) * 2^(-2* 7) )   n =  7   d_n = 0 
assign u[4'b0000] [07] = 21'h 000000;  // +0.0000000000000000 = 2^ 8 * ln( 1 +  0 * 2^(- 8+1) + ( 0^2+ 0^2) * 2^(-2* 8) )   n =  8   d_n = 0 
assign u[4'b0000] [08] = 21'h 000000;  // +0.0000000000000000 = 2^ 9 * ln( 1 +  0 * 2^(- 9+1) + ( 0^2+ 0^2) * 2^(-2* 9) )   n =  9   d_n = 0 
assign u[4'b0000] [09] = 21'h 000000;  // +0.0000000000000000 = 2^10 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = 0 
assign u[4'b0000] [10] = 21'h 000000;  // +0.0000000000000000 = 2^11 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = 0 
assign u[4'b0000] [11] = 21'h 000000;  // +0.0000000000000000 = 2^12 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = 0 
assign u[4'b0000] [12] = 21'h 000000;  // +0.0000000000000000 = 2^13 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = 0 
assign u[4'b0000] [13] = 21'h 000000;  // +0.0000000000000000 = 2^14 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = 0 
assign u[4'b0000] [14] = 21'h 000000;  // +0.0000000000000000 = 2^15 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = 0 
assign u[4'b0000] [15] = 21'h 000000;  // +0.0000000000000000 = 2^16 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = 0 
assign u[4'b0000] [16] = 21'h 000000;  // +0.0000000000000000 = 2^17 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = 0 
assign u[4'b0000] [17] = 21'h 000000;  // +0.0000000000000000 = 2^18 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = 0 
assign u[4'b0000] [18] = 21'h 000000;  // +0.0000000000000000 = 2^19 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = 0 
assign u[4'b0000] [19] = 21'h 000000;  // +0.0000000000000000 = 2^20 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = 0 
assign u[4'b0000] [20] = 21'h 000000;  // +0.0000000000000000 = 2^21 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = 0 
assign u[4'b0000] [21] = 21'h 000000;  // +0.0000000000000000 = 2^22 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = 0 
assign u[4'b0000] [22] = 21'h 000000;  // +0.0000000000000000 = 2^23 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = 0 
assign u[4'b0000] [23] = 21'h 000000;  // +0.0000000000000000 = 2^24 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = 0 
assign u[4'b0000] [24] = 21'h 000000;  // +0.0000000000000000 = 2^25 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = 0 
assign u[4'b0000] [25] = 21'h 000000;  // +0.0000000000000000 = 2^26 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = 0 
assign u[4'b0000] [26] = 21'h 000000;  // +0.0000000000000000 = 2^27 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = 0 
assign u[4'b0000] [27] = 21'h 000000;  // +0.0000000000000000 = 2^28 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = 0 
assign u[4'b0000] [28] = 21'h 000000;  // +0.0000000000000000 = 2^29 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = 0 
assign u[4'b0000] [29] = 21'h 000000;  // +0.0000000000000000 = 2^30 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = 0 
assign u[4'b0000] [30] = 21'h 000000;  // +0.0000000000000000 = 2^31 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = 0 
assign u[4'b0000] [31] = 21'h 000000;  // +0.0000000000000000 = 2^32 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = 0 
assign u[4'b0000] [32] = 21'h 000000;  // +0.0000000000000000 = 2^33 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = 0 
assign u[4'b0000] [33] = 21'h 000000;  // +0.0000000000000000 = 2^34 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = 0 
assign u[4'b0000] [34] = 21'h 000000;  // +0.0000000000000000 = 2^35 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = 0 
assign u[4'b0000] [35] = 21'h 000000;  // +0.0000000000000000 = 2^36 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = 0 
assign u[4'b0000] [36] = 21'h 000000;  // +0.0000000000000000 = 2^37 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = 0 
assign u[4'b0000] [37] = 21'h 000000;  // +0.0000000000000000 = 2^38 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = 0 
assign u[4'b0000] [38] = 21'h 000000;  // +0.0000000000000000 = 2^39 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = 0 
assign u[4'b0000] [39] = 21'h 000000;  // +0.0000000000000000 = 2^40 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = 0 
assign u[4'b0000] [40] = 21'h 000000;  // +0.0000000000000000 = 2^41 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = 0 
assign u[4'b0000] [41] = 21'h 000000;  // +0.0000000000000000 = 2^42 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = 0 
assign u[4'b0000] [42] = 21'h 000000;  // +0.0000000000000000 = 2^43 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = 0 
assign u[4'b0000] [43] = 21'h 000000;  // +0.0000000000000000 = 2^44 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = 0 
assign u[4'b0000] [44] = 21'h 000000;  // +0.0000000000000000 = 2^45 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = 0 
assign u[4'b0000] [45] = 21'h 000000;  // +0.0000000000000000 = 2^46 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = 0 
assign u[4'b0000] [46] = 21'h 000000;  // +0.0000000000000000 = 2^47 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = 0 
assign u[4'b0000] [47] = 21'h 000000;  // +0.0000000000000000 = 2^48 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = 0 
assign u[4'b0000] [48] = 21'h 000000;  // +0.0000000000000000 = 2^49 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = 0 
assign u[4'b0000] [49] = 21'h 000000;  // +0.0000000000000000 = 2^50 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = 0 
assign u[4'b0000] [50] = 21'h 000000;  // +0.0000000000000000 = 2^51 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = 0 
assign u[4'b0000] [51] = 21'h 000000;  // +0.0000000000000000 = 2^52 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = 0 
assign u[4'b0000] [52] = 21'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = 0 
assign u[4'b0000] [53] = 21'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = 0 
assign u[4'b0000] [54] = 21'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = 0 
assign u[4'b0000] [55] = 21'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = 0 
assign u[4'b0000] [56] = 21'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = 0 
assign u[4'b0000] [57] = 21'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = 0 
assign u[4'b0000] [58] = 21'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = 0 
assign u[4'b0000] [59] = 21'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = 0 
assign u[4'b0000] [60] = 21'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = 0 
assign u[4'b0000] [61] = 21'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = 0 
assign u[4'b0000] [62] = 21'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = 0 
assign u[4'b0000] [63] = 21'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = 0 
assign u[4'b0001] [00] = 21'h 00067C;  // +1.6218604324326575 = 2^ 1 * ln( 1 +  1 * 2^(- 1+1) + ( 1^2+ 0^2) * 2^(-2* 1) )   n =  1   d_n = 1 
assign u[4'b0001] [01] = 21'h 000723;  // +1.7851484105136781 = 2^ 2 * ln( 1 +  1 * 2^(- 2+1) + ( 1^2+ 0^2) * 2^(-2* 2) )   n =  2   d_n = 1 
assign u[4'b0001] [02] = 21'h 000789;  // +1.8845285705021353 = 2^ 3 * ln( 1 +  1 * 2^(- 3+1) + ( 1^2+ 0^2) * 2^(-2* 3) )   n =  3   d_n = 1 
assign u[4'b0001] [03] = 21'h 0007C2;  // +1.9399878981259149 = 2^ 4 * ln( 1 +  1 * 2^(- 4+1) + ( 1^2+ 0^2) * 2^(-2* 4) )   n =  4   d_n = 1 
assign u[4'b0001] [04] = 21'h 0007E0;  // +1.9693861546722360 = 2^ 5 * ln( 1 +  1 * 2^(- 5+1) + ( 1^2+ 0^2) * 2^(-2* 5) )   n =  5   d_n = 1 
assign u[4'b0001] [05] = 21'h 0007F0;  // +1.9845358766035526 = 2^ 6 * ln( 1 +  1 * 2^(- 6+1) + ( 1^2+ 0^2) * 2^(-2* 6) )   n =  6   d_n = 1 
assign u[4'b0001] [06] = 21'h 0007F8;  // +1.9922279531660669 = 2^ 7 * ln( 1 +  1 * 2^(- 7+1) + ( 1^2+ 0^2) * 2^(-2* 7) )   n =  7   d_n = 1 
assign u[4'b0001] [07] = 21'h 0007FC;  // +1.9961038928165493 = 2^ 8 * ln( 1 +  1 * 2^(- 8+1) + ( 1^2+ 0^2) * 2^(-2* 8) )   n =  8   d_n = 1 
assign u[4'b0001] [08] = 21'h 0007FE;  // +1.9980494144120313 = 2^ 9 * ln( 1 +  1 * 2^(- 9+1) + ( 1^2+ 0^2) * 2^(-2* 9) )   n =  9   d_n = 1 
assign u[4'b0001] [09] = 21'h 0007FF;  // +1.9990240728175799 = 2^10 * ln( 1 +  1 * 2^(-10+1) + ( 1^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = 1 
assign u[4'b0001] [10] = 21'h 0007FF;  // +1.9995118776375345 = 2^11 * ln( 1 +  1 * 2^(-11+1) + ( 1^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = 1 
assign u[4'b0001] [11] = 21'h 0007FF;  // +1.9997558991041553 = 2^12 * ln( 1 +  1 * 2^(-12+1) + ( 1^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = 1 
assign u[4'b0001] [12] = 21'h 0007FF;  // +1.9998779396206980 = 2^13 * ln( 1 +  1 * 2^(-13+1) + ( 1^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = 1 
assign u[4'b0001] [13] = 21'h 0007FF;  // +1.9999389673271633 = 2^14 * ln( 1 +  1 * 2^(-14+1) + ( 1^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = 1 
assign u[4'b0001] [14] = 21'h 0007FF;  // +1.9999694830427426 = 2^15 * ln( 1 +  1 * 2^(-15+1) + ( 1^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = 1 
assign u[4'b0001] [15] = 21'h 0007FF;  // +1.9999847413661562 = 2^16 * ln( 1 +  1 * 2^(-16+1) + ( 1^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = 1 
assign u[4'b0001] [16] = 21'h 0007FF;  // +1.9999923706442737 = 2^17 * ln( 1 +  1 * 2^(-17+1) + ( 1^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = 1 
assign u[4'b0001] [17] = 21'h 0007FF;  // +1.9999961853124357 = 2^18 * ln( 1 +  1 * 2^(-18+1) + ( 1^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = 1 
assign u[4'b0001] [18] = 21'h 0007FF;  // +1.9999980926537926 = 2^19 * ln( 1 +  1 * 2^(-19+1) + ( 1^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = 1 
assign u[4'b0001] [19] = 21'h 0007FF;  // +1.9999990463262900 = 2^20 * ln( 1 +  1 * 2^(-20+1) + ( 1^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = 1 
assign u[4'b0001] [20] = 21'h 0007FF;  // +1.9999995231629935 = 2^21 * ln( 1 +  1 * 2^(-21+1) + ( 1^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = 1 
assign u[4'b0001] [21] = 21'h 0007FF;  // +1.9999997615814589 = 2^22 * ln( 1 +  1 * 2^(-22+1) + ( 1^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = 1 
assign u[4'b0001] [22] = 21'h 0007FF;  // +1.9999998807907200 = 2^23 * ln( 1 +  1 * 2^(-23+1) + ( 1^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = 1 
assign u[4'b0001] [23] = 21'h 0007FF;  // +1.9999999403953577 = 2^24 * ln( 1 +  1 * 2^(-24+1) + ( 1^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = 1 
assign u[4'b0001] [24] = 21'h 0007FF;  // +1.9999999701976783 = 2^25 * ln( 1 +  1 * 2^(-25+1) + ( 1^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = 1 
assign u[4'b0001] [25] = 21'h 0007FF;  // +1.9999999850988390 = 2^26 * ln( 1 +  1 * 2^(-26+1) + ( 1^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = 1 
assign u[4'b0001] [26] = 21'h 0007FF;  // +1.9999999925494194 = 2^27 * ln( 1 +  1 * 2^(-27+1) + ( 1^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = 1 
assign u[4'b0001] [27] = 21'h 0007FF;  // +1.9999999962747097 = 2^28 * ln( 1 +  1 * 2^(-28+1) + ( 1^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = 1 
assign u[4'b0001] [28] = 21'h 0007FF;  // +1.9999999981373549 = 2^29 * ln( 1 +  1 * 2^(-29+1) + ( 1^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = 1 
assign u[4'b0001] [29] = 21'h 0007FF;  // +1.9999999990686774 = 2^30 * ln( 1 +  1 * 2^(-30+1) + ( 1^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = 1 
assign u[4'b0001] [30] = 21'h 0007FF;  // +1.9999999995343387 = 2^31 * ln( 1 +  1 * 2^(-31+1) + ( 1^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = 1 
assign u[4'b0001] [31] = 21'h 0007FF;  // +1.9999999997671694 = 2^32 * ln( 1 +  1 * 2^(-32+1) + ( 1^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = 1 
assign u[4'b0001] [32] = 21'h 0007FF;  // +1.9999999998835847 = 2^33 * ln( 1 +  1 * 2^(-33+1) + ( 1^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = 1 
assign u[4'b0001] [33] = 21'h 0007FF;  // +1.9999999999417923 = 2^34 * ln( 1 +  1 * 2^(-34+1) + ( 1^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = 1 
assign u[4'b0001] [34] = 21'h 0007FF;  // +1.9999999999708962 = 2^35 * ln( 1 +  1 * 2^(-35+1) + ( 1^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = 1 
assign u[4'b0001] [35] = 21'h 0007FF;  // +1.9999999999854481 = 2^36 * ln( 1 +  1 * 2^(-36+1) + ( 1^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = 1 
assign u[4'b0001] [36] = 21'h 0007FF;  // +1.9999999999927240 = 2^37 * ln( 1 +  1 * 2^(-37+1) + ( 1^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = 1 
assign u[4'b0001] [37] = 21'h 0007FF;  // +1.9999999999963620 = 2^38 * ln( 1 +  1 * 2^(-38+1) + ( 1^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = 1 
assign u[4'b0001] [38] = 21'h 0007FF;  // +1.9999999999981810 = 2^39 * ln( 1 +  1 * 2^(-39+1) + ( 1^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = 1 
assign u[4'b0001] [39] = 21'h 0007FF;  // +1.9999999999990905 = 2^40 * ln( 1 +  1 * 2^(-40+1) + ( 1^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = 1 
assign u[4'b0001] [40] = 21'h 0007FF;  // +1.9999999999995453 = 2^41 * ln( 1 +  1 * 2^(-41+1) + ( 1^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = 1 
assign u[4'b0001] [41] = 21'h 0007FF;  // +1.9999999999997726 = 2^42 * ln( 1 +  1 * 2^(-42+1) + ( 1^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = 1 
assign u[4'b0001] [42] = 21'h 0007FF;  // +1.9999999999998863 = 2^43 * ln( 1 +  1 * 2^(-43+1) + ( 1^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = 1 
assign u[4'b0001] [43] = 21'h 0007FF;  // +1.9999999999999432 = 2^44 * ln( 1 +  1 * 2^(-44+1) + ( 1^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = 1 
assign u[4'b0001] [44] = 21'h 0007FF;  // +1.9999999999999716 = 2^45 * ln( 1 +  1 * 2^(-45+1) + ( 1^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = 1 
assign u[4'b0001] [45] = 21'h 0007FF;  // +1.9999999999999858 = 2^46 * ln( 1 +  1 * 2^(-46+1) + ( 1^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = 1 
assign u[4'b0001] [46] = 21'h 0007FF;  // +1.9999999999999929 = 2^47 * ln( 1 +  1 * 2^(-47+1) + ( 1^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = 1 
assign u[4'b0001] [47] = 21'h 0007FF;  // +1.9999999999999964 = 2^48 * ln( 1 +  1 * 2^(-48+1) + ( 1^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = 1 
assign u[4'b0001] [48] = 21'h 0007FF;  // +1.9999999999999982 = 2^49 * ln( 1 +  1 * 2^(-49+1) + ( 1^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = 1 
assign u[4'b0001] [49] = 21'h 0007FF;  // +1.9999999999999991 = 2^50 * ln( 1 +  1 * 2^(-50+1) + ( 1^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = 1 
assign u[4'b0001] [50] = 21'h 0007FF;  // +1.9999999999999996 = 2^51 * ln( 1 +  1 * 2^(-51+1) + ( 1^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = 1 
assign u[4'b0001] [51] = 21'h 0007FF;  // +1.9999999999999998 = 2^52 * ln( 1 +  1 * 2^(-52+1) + ( 1^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = 1 
assign u[4'b0001] [52] = 21'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  1 * 2^(-53+1) + ( 1^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = 1 
assign u[4'b0001] [53] = 21'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  1 * 2^(-54+1) + ( 1^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = 1 
assign u[4'b0001] [54] = 21'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  1 * 2^(-55+1) + ( 1^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = 1 
assign u[4'b0001] [55] = 21'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  1 * 2^(-56+1) + ( 1^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = 1 
assign u[4'b0001] [56] = 21'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  1 * 2^(-57+1) + ( 1^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = 1 
assign u[4'b0001] [57] = 21'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  1 * 2^(-58+1) + ( 1^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = 1 
assign u[4'b0001] [58] = 21'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  1 * 2^(-59+1) + ( 1^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = 1 
assign u[4'b0001] [59] = 21'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  1 * 2^(-60+1) + ( 1^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = 1 
assign u[4'b0001] [60] = 21'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  1 * 2^(-61+1) + ( 1^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = 1 
assign u[4'b0001] [61] = 21'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  1 * 2^(-62+1) + ( 1^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = 1 
assign u[4'b0001] [62] = 21'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  1 * 2^(-63+1) + ( 1^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = 1 
assign u[4'b0001] [63] = 21'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  1 * 2^(-64+1) + ( 1^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = 1 
assign u[4'b0010] [00] = 21'h 000000;  // +0.0000000000000000 = 2^ 1 * ln( 1 +  0 * 2^(- 1+1) + ( 0^2+ 0^2) * 2^(-2* 1) )   n =  1   d_n = -0 
assign u[4'b0010] [01] = 21'h 000000;  // +0.0000000000000000 = 2^ 2 * ln( 1 +  0 * 2^(- 2+1) + ( 0^2+ 0^2) * 2^(-2* 2) )   n =  2   d_n = -0 
assign u[4'b0010] [02] = 21'h 000000;  // +0.0000000000000000 = 2^ 3 * ln( 1 +  0 * 2^(- 3+1) + ( 0^2+ 0^2) * 2^(-2* 3) )   n =  3   d_n = -0 
assign u[4'b0010] [03] = 21'h 000000;  // +0.0000000000000000 = 2^ 4 * ln( 1 +  0 * 2^(- 4+1) + ( 0^2+ 0^2) * 2^(-2* 4) )   n =  4   d_n = -0 
assign u[4'b0010] [04] = 21'h 000000;  // +0.0000000000000000 = 2^ 5 * ln( 1 +  0 * 2^(- 5+1) + ( 0^2+ 0^2) * 2^(-2* 5) )   n =  5   d_n = -0 
assign u[4'b0010] [05] = 21'h 000000;  // +0.0000000000000000 = 2^ 6 * ln( 1 +  0 * 2^(- 6+1) + ( 0^2+ 0^2) * 2^(-2* 6) )   n =  6   d_n = -0 
assign u[4'b0010] [06] = 21'h 000000;  // +0.0000000000000000 = 2^ 7 * ln( 1 +  0 * 2^(- 7+1) + ( 0^2+ 0^2) * 2^(-2* 7) )   n =  7   d_n = -0 
assign u[4'b0010] [07] = 21'h 000000;  // +0.0000000000000000 = 2^ 8 * ln( 1 +  0 * 2^(- 8+1) + ( 0^2+ 0^2) * 2^(-2* 8) )   n =  8   d_n = -0 
assign u[4'b0010] [08] = 21'h 000000;  // +0.0000000000000000 = 2^ 9 * ln( 1 +  0 * 2^(- 9+1) + ( 0^2+ 0^2) * 2^(-2* 9) )   n =  9   d_n = -0 
assign u[4'b0010] [09] = 21'h 000000;  // +0.0000000000000000 = 2^10 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = -0 
assign u[4'b0010] [10] = 21'h 000000;  // +0.0000000000000000 = 2^11 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = -0 
assign u[4'b0010] [11] = 21'h 000000;  // +0.0000000000000000 = 2^12 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = -0 
assign u[4'b0010] [12] = 21'h 000000;  // +0.0000000000000000 = 2^13 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = -0 
assign u[4'b0010] [13] = 21'h 000000;  // +0.0000000000000000 = 2^14 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = -0 
assign u[4'b0010] [14] = 21'h 000000;  // +0.0000000000000000 = 2^15 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = -0 
assign u[4'b0010] [15] = 21'h 000000;  // +0.0000000000000000 = 2^16 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = -0 
assign u[4'b0010] [16] = 21'h 000000;  // +0.0000000000000000 = 2^17 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = -0 
assign u[4'b0010] [17] = 21'h 000000;  // +0.0000000000000000 = 2^18 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = -0 
assign u[4'b0010] [18] = 21'h 000000;  // +0.0000000000000000 = 2^19 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = -0 
assign u[4'b0010] [19] = 21'h 000000;  // +0.0000000000000000 = 2^20 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = -0 
assign u[4'b0010] [20] = 21'h 000000;  // +0.0000000000000000 = 2^21 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = -0 
assign u[4'b0010] [21] = 21'h 000000;  // +0.0000000000000000 = 2^22 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = -0 
assign u[4'b0010] [22] = 21'h 000000;  // +0.0000000000000000 = 2^23 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = -0 
assign u[4'b0010] [23] = 21'h 000000;  // +0.0000000000000000 = 2^24 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = -0 
assign u[4'b0010] [24] = 21'h 000000;  // +0.0000000000000000 = 2^25 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = -0 
assign u[4'b0010] [25] = 21'h 000000;  // +0.0000000000000000 = 2^26 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = -0 
assign u[4'b0010] [26] = 21'h 000000;  // +0.0000000000000000 = 2^27 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = -0 
assign u[4'b0010] [27] = 21'h 000000;  // +0.0000000000000000 = 2^28 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = -0 
assign u[4'b0010] [28] = 21'h 000000;  // +0.0000000000000000 = 2^29 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = -0 
assign u[4'b0010] [29] = 21'h 000000;  // +0.0000000000000000 = 2^30 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = -0 
assign u[4'b0010] [30] = 21'h 000000;  // +0.0000000000000000 = 2^31 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = -0 
assign u[4'b0010] [31] = 21'h 000000;  // +0.0000000000000000 = 2^32 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = -0 
assign u[4'b0010] [32] = 21'h 000000;  // +0.0000000000000000 = 2^33 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = -0 
assign u[4'b0010] [33] = 21'h 000000;  // +0.0000000000000000 = 2^34 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = -0 
assign u[4'b0010] [34] = 21'h 000000;  // +0.0000000000000000 = 2^35 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = -0 
assign u[4'b0010] [35] = 21'h 000000;  // +0.0000000000000000 = 2^36 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = -0 
assign u[4'b0010] [36] = 21'h 000000;  // +0.0000000000000000 = 2^37 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = -0 
assign u[4'b0010] [37] = 21'h 000000;  // +0.0000000000000000 = 2^38 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = -0 
assign u[4'b0010] [38] = 21'h 000000;  // +0.0000000000000000 = 2^39 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = -0 
assign u[4'b0010] [39] = 21'h 000000;  // +0.0000000000000000 = 2^40 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = -0 
assign u[4'b0010] [40] = 21'h 000000;  // +0.0000000000000000 = 2^41 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = -0 
assign u[4'b0010] [41] = 21'h 000000;  // +0.0000000000000000 = 2^42 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = -0 
assign u[4'b0010] [42] = 21'h 000000;  // +0.0000000000000000 = 2^43 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = -0 
assign u[4'b0010] [43] = 21'h 000000;  // +0.0000000000000000 = 2^44 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = -0 
assign u[4'b0010] [44] = 21'h 000000;  // +0.0000000000000000 = 2^45 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = -0 
assign u[4'b0010] [45] = 21'h 000000;  // +0.0000000000000000 = 2^46 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = -0 
assign u[4'b0010] [46] = 21'h 000000;  // +0.0000000000000000 = 2^47 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = -0 
assign u[4'b0010] [47] = 21'h 000000;  // +0.0000000000000000 = 2^48 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = -0 
assign u[4'b0010] [48] = 21'h 000000;  // +0.0000000000000000 = 2^49 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = -0 
assign u[4'b0010] [49] = 21'h 000000;  // +0.0000000000000000 = 2^50 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = -0 
assign u[4'b0010] [50] = 21'h 000000;  // +0.0000000000000000 = 2^51 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = -0 
assign u[4'b0010] [51] = 21'h 000000;  // +0.0000000000000000 = 2^52 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = -0 
assign u[4'b0010] [52] = 21'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = -0 
assign u[4'b0010] [53] = 21'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = -0 
assign u[4'b0010] [54] = 21'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = -0 
assign u[4'b0010] [55] = 21'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = -0 
assign u[4'b0010] [56] = 21'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = -0 
assign u[4'b0010] [57] = 21'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = -0 
assign u[4'b0010] [58] = 21'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = -0 
assign u[4'b0010] [59] = 21'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = -0 
assign u[4'b0010] [60] = 21'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = -0 
assign u[4'b0010] [61] = 21'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = -0 
assign u[4'b0010] [62] = 21'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = -0 
assign u[4'b0010] [63] = 21'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = -0 
assign u[4'b0011] [00] = 21'h 1FF4E8;  // -2.7725887222397811 = 2^ 1 * ln( 1 + -1 * 2^(- 1+1) + (-1^2+ 0^2) * 2^(-2* 1) )   n =  1   d_n = -1 
assign u[4'b0011] [01] = 21'h 1FF6CB;  // -2.3014565796142472 = 2^ 2 * ln( 1 + -1 * 2^(- 2+1) + (-1^2+ 0^2) * 2^(-2* 2) )   n =  2   d_n = -1 
assign u[4'b0011] [02] = 21'h 1FF774;  // -2.1365022819923620 = 2^ 3 * ln( 1 + -1 * 2^(- 3+1) + (-1^2+ 0^2) * 2^(-2* 3) )   n =  3   d_n = -1 
assign u[4'b0011] [03] = 21'h 1FF7BD;  // -2.0652326764022777 = 2^ 4 * ln( 1 + -1 * 2^(- 4+1) + (-1^2+ 0^2) * 2^(-2* 4) )   n =  4   d_n = -1 
assign u[4'b0011] [04] = 21'h 1FF7DF;  // -2.0319166921331391 = 2^ 5 * ln( 1 + -1 * 2^(- 5+1) + (-1^2+ 0^2) * 2^(-2* 5) )   n =  5   d_n = -1 
assign u[4'b0011] [05] = 21'h 1FF7EF;  // -2.0157896919218135 = 2^ 6 * ln( 1 + -1 * 2^(- 6+1) + (-1^2+ 0^2) * 2^(-2* 6) )   n =  6   d_n = -1 
assign u[4'b0011] [06] = 21'h 1FF7F7;  // -2.0078534300226285 = 2^ 7 * ln( 1 + -1 * 2^(- 7+1) + (-1^2+ 0^2) * 2^(-2* 7) )   n =  7   d_n = -1 
assign u[4'b0011] [07] = 21'h 1FF7FB;  // -2.0039164524218003 = 2^ 8 * ln( 1 + -1 * 2^(- 8+1) + (-1^2+ 0^2) * 2^(-2* 8) )   n =  8   d_n = -1 
assign u[4'b0011] [08] = 21'h 1FF7FD;  // -2.0019556718626310 = 2^ 9 * ln( 1 + -1 * 2^(- 9+1) + (-1^2+ 0^2) * 2^(-2* 9) )   n =  9   d_n = -1 
assign u[4'b0011] [09] = 21'h 1FF7FE;  // -2.0009771987489029 = 2^10 * ln( 1 + -1 * 2^(-10+1) + (-1^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = -1 
assign u[4'b0011] [10] = 21'h 1FF7FF;  // -2.0004884402539500 = 2^11 * ln( 1 + -1 * 2^(-11+1) + (-1^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = -1 
assign u[4'b0011] [11] = 21'h 1FF7FF;  // -2.0002441803687074 = 2^12 * ln( 1 + -1 * 2^(-12+1) + (-1^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = -1 
assign u[4'b0011] [12] = 21'h 1FF7FF;  // -2.0001220802475173 = 2^13 * ln( 1 + -1 * 2^(-13+1) + (-1^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = -1 
assign u[4'b0011] [13] = 21'h 1FF7FF;  // -2.0000610376398904 = 2^14 * ln( 1 + -1 * 2^(-14+1) + (-1^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = -1 
assign u[4'b0011] [14] = 21'h 1FF7FF;  // -2.0000305181990208 = 2^15 * ln( 1 + -1 * 2^(-15+1) + (-1^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = -1 
assign u[4'b0011] [15] = 21'h 1FF7FF;  // -2.0000152589442846 = 2^16 * ln( 1 + -1 * 2^(-16+1) + (-1^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = -1 
assign u[4'b0011] [16] = 21'h 1FF7FF;  // -2.0000076294333367 = 2^17 * ln( 1 + -1 * 2^(-17+1) + (-1^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = -1 
assign u[4'b0011] [17] = 21'h 1FF7FF;  // -2.0000038147069668 = 2^18 * ln( 1 + -1 * 2^(-18+1) + (-1^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = -1 
assign u[4'b0011] [18] = 21'h 1FF7FF;  // -2.0000019073510580 = 2^19 * ln( 1 + -1 * 2^(-19+1) + (-1^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = -1 
assign u[4'b0011] [19] = 21'h 1FF7FF;  // -2.0000009536749226 = 2^20 * ln( 1 + -1 * 2^(-20+1) + (-1^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = -1 
assign u[4'b0011] [20] = 21'h 1FF7FF;  // -2.0000004768373096 = 2^21 * ln( 1 + -1 * 2^(-21+1) + (-1^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = -1 
assign u[4'b0011] [21] = 21'h 1FF7FF;  // -2.0000002384186168 = 2^22 * ln( 1 + -1 * 2^(-22+1) + (-1^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = -1 
assign u[4'b0011] [22] = 21'h 1FF7FF;  // -2.0000001192092989 = 2^23 * ln( 1 + -1 * 2^(-23+1) + (-1^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = -1 
assign u[4'b0011] [23] = 21'h 1FF7FF;  // -2.0000000596046470 = 2^24 * ln( 1 + -1 * 2^(-24+1) + (-1^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = -1 
assign u[4'b0011] [24] = 21'h 1FF7FF;  // -2.0000000298023228 = 2^25 * ln( 1 + -1 * 2^(-25+1) + (-1^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = -1 
assign u[4'b0011] [25] = 21'h 1FF7FF;  // -2.0000000149011612 = 2^26 * ln( 1 + -1 * 2^(-26+1) + (-1^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = -1 
assign u[4'b0011] [26] = 21'h 1FF7FF;  // -2.0000000074505806 = 2^27 * ln( 1 + -1 * 2^(-27+1) + (-1^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = -1 
assign u[4'b0011] [27] = 21'h 1FF7FF;  // -2.0000000037252903 = 2^28 * ln( 1 + -1 * 2^(-28+1) + (-1^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = -1 
assign u[4'b0011] [28] = 21'h 1FF7FF;  // -2.0000000018626451 = 2^29 * ln( 1 + -1 * 2^(-29+1) + (-1^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = -1 
assign u[4'b0011] [29] = 21'h 1FF7FF;  // -2.0000000009313226 = 2^30 * ln( 1 + -1 * 2^(-30+1) + (-1^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = -1 
assign u[4'b0011] [30] = 21'h 1FF7FF;  // -2.0000000004656613 = 2^31 * ln( 1 + -1 * 2^(-31+1) + (-1^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = -1 
assign u[4'b0011] [31] = 21'h 1FF7FF;  // -2.0000000002328306 = 2^32 * ln( 1 + -1 * 2^(-32+1) + (-1^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = -1 
assign u[4'b0011] [32] = 21'h 1FF7FF;  // -2.0000000001164153 = 2^33 * ln( 1 + -1 * 2^(-33+1) + (-1^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = -1 
assign u[4'b0011] [33] = 21'h 1FF7FF;  // -2.0000000000582077 = 2^34 * ln( 1 + -1 * 2^(-34+1) + (-1^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = -1 
assign u[4'b0011] [34] = 21'h 1FF7FF;  // -2.0000000000291038 = 2^35 * ln( 1 + -1 * 2^(-35+1) + (-1^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = -1 
assign u[4'b0011] [35] = 21'h 1FF7FF;  // -2.0000000000145519 = 2^36 * ln( 1 + -1 * 2^(-36+1) + (-1^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = -1 
assign u[4'b0011] [36] = 21'h 1FF7FF;  // -2.0000000000072760 = 2^37 * ln( 1 + -1 * 2^(-37+1) + (-1^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = -1 
assign u[4'b0011] [37] = 21'h 1FF7FF;  // -2.0000000000036380 = 2^38 * ln( 1 + -1 * 2^(-38+1) + (-1^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = -1 
assign u[4'b0011] [38] = 21'h 1FF7FF;  // -2.0000000000018190 = 2^39 * ln( 1 + -1 * 2^(-39+1) + (-1^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = -1 
assign u[4'b0011] [39] = 21'h 1FF7FF;  // -2.0000000000009095 = 2^40 * ln( 1 + -1 * 2^(-40+1) + (-1^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = -1 
assign u[4'b0011] [40] = 21'h 1FF7FF;  // -2.0000000000004547 = 2^41 * ln( 1 + -1 * 2^(-41+1) + (-1^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = -1 
assign u[4'b0011] [41] = 21'h 1FF7FF;  // -2.0000000000002274 = 2^42 * ln( 1 + -1 * 2^(-42+1) + (-1^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = -1 
assign u[4'b0011] [42] = 21'h 1FF800;  // -2.0000000000001137 = 2^43 * ln( 1 + -1 * 2^(-43+1) + (-1^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = -1 
assign u[4'b0011] [43] = 21'h 1FF800;  // -2.0000000000000568 = 2^44 * ln( 1 + -1 * 2^(-44+1) + (-1^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = -1 
assign u[4'b0011] [44] = 21'h 1FF800;  // -2.0000000000000284 = 2^45 * ln( 1 + -1 * 2^(-45+1) + (-1^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = -1 
assign u[4'b0011] [45] = 21'h 1FF800;  // -2.0000000000000142 = 2^46 * ln( 1 + -1 * 2^(-46+1) + (-1^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = -1 
assign u[4'b0011] [46] = 21'h 1FF800;  // -2.0000000000000071 = 2^47 * ln( 1 + -1 * 2^(-47+1) + (-1^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = -1 
assign u[4'b0011] [47] = 21'h 1FF800;  // -2.0000000000000036 = 2^48 * ln( 1 + -1 * 2^(-48+1) + (-1^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = -1 
assign u[4'b0011] [48] = 21'h 1FF800;  // -2.0000000000000018 = 2^49 * ln( 1 + -1 * 2^(-49+1) + (-1^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = -1 
assign u[4'b0011] [49] = 21'h 1FF800;  // -2.0000000000000009 = 2^50 * ln( 1 + -1 * 2^(-50+1) + (-1^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = -1 
assign u[4'b0011] [50] = 21'h 1FF800;  // -2.0000000000000004 = 2^51 * ln( 1 + -1 * 2^(-51+1) + (-1^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = -1 
assign u[4'b0011] [51] = 21'h 1FF800;  // -2.0000000000000004 = 2^52 * ln( 1 + -1 * 2^(-52+1) + (-1^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = -1 
assign u[4'b0011] [52] = 21'h 1FF800;  // -2.0000000000000000 = 2^53 * ln( 1 + -1 * 2^(-53+1) + (-1^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = -1 
assign u[4'b0011] [53] = 21'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 + -1 * 2^(-54+1) + (-1^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = -1 
assign u[4'b0011] [54] = 21'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 + -1 * 2^(-55+1) + (-1^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = -1 
assign u[4'b0011] [55] = 21'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 + -1 * 2^(-56+1) + (-1^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = -1 
assign u[4'b0011] [56] = 21'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 + -1 * 2^(-57+1) + (-1^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = -1 
assign u[4'b0011] [57] = 21'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 + -1 * 2^(-58+1) + (-1^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = -1 
assign u[4'b0011] [58] = 21'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 + -1 * 2^(-59+1) + (-1^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = -1 
assign u[4'b0011] [59] = 21'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 + -1 * 2^(-60+1) + (-1^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = -1 
assign u[4'b0011] [60] = 21'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 + -1 * 2^(-61+1) + (-1^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = -1 
assign u[4'b0011] [61] = 21'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 + -1 * 2^(-62+1) + (-1^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = -1 
assign u[4'b0011] [62] = 21'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 + -1 * 2^(-63+1) + (-1^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = -1 
assign u[4'b0011] [63] = 21'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 + -1 * 2^(-64+1) + (-1^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = -1 
assign u[4'b0100] [00] = 21'h 0001C8;  // +0.4462871026284197 = 2^ 1 * ln( 1 +  0 * 2^(- 1+1) + ( 0^2+ 1^2) * 2^(-2* 1) )   n =  1   d_n = 0+1i 
assign u[4'b0100] [01] = 21'h 0000F8;  // +0.2424984872657394 = 2^ 2 * ln( 1 +  0 * 2^(- 2+1) + ( 0^2+ 1^2) * 2^(-2* 2) )   n =  2   d_n = 0+1i 
assign u[4'b0100] [02] = 21'h 00007F;  // +0.1240334922877210 = 2^ 3 * ln( 1 +  0 * 2^(- 3+1) + ( 0^2+ 1^2) * 2^(-2* 3) )   n =  3   d_n = 0+1i 
assign u[4'b0100] [03] = 21'h 00003F;  // +0.0623782466505195 = 2^ 4 * ln( 1 +  0 * 2^(- 4+1) + ( 0^2+ 1^2) * 2^(-2* 4) )   n =  4   d_n = 0+1i 
assign u[4'b0100] [04] = 21'h 00001F;  // +0.0312347511377731 = 2^ 5 * ln( 1 +  0 * 2^(- 5+1) + ( 0^2+ 1^2) * 2^(-2* 5) )   n =  5   d_n = 0+1i 
assign u[4'b0100] [05] = 21'h 00000F;  // +0.0156230929617406 = 2^ 6 * ln( 1 +  0 * 2^(- 6+1) + ( 0^2+ 1^2) * 2^(-2* 6) )   n =  6   d_n = 0+1i 
assign u[4'b0100] [06] = 21'h 000007;  // +0.0078122615911219 = 2^ 7 * ln( 1 +  0 * 2^(- 7+1) + ( 0^2+ 1^2) * 2^(-2* 7) )   n =  7   d_n = 0+1i 
assign u[4'b0100] [07] = 21'h 000003;  // +0.0039062201979808 = 2^ 8 * ln( 1 +  0 * 2^(- 8+1) + ( 0^2+ 1^2) * 2^(-2* 8) )   n =  8   d_n = 0+1i 
assign u[4'b0100] [08] = 21'h 000001;  // +0.0019531212747156 = 2^ 9 * ln( 1 +  0 * 2^(- 9+1) + ( 0^2+ 1^2) * 2^(-2* 9) )   n =  9   d_n = 0+1i 
assign u[4'b0100] [09] = 21'h 000000;  // +0.0009765620343389 = 2^10 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 1^2) * 2^(-2*10) )   n = 10   d_n = 0+1i 
assign u[4'b0100] [10] = 21'h 000000;  // +0.0004882811917923 = 2^11 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 1^2) * 2^(-2*11) )   n = 11   d_n = 0+1i 
assign u[4'b0100] [11] = 21'h 000000;  // +0.0002441406177240 = 2^12 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 1^2) * 2^(-2*12) )   n = 12   d_n = 0+1i 
assign u[4'b0100] [12] = 21'h 000000;  // +0.0001220703120453 = 2^13 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 1^2) * 2^(-2*13) )   n = 13   d_n = 0+1i 
assign u[4'b0100] [13] = 21'h 000000;  // +0.0000610351561932 = 2^14 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 1^2) * 2^(-2*14) )   n = 14   d_n = 0+1i 
assign u[4'b0100] [14] = 21'h 000000;  // +0.0000305175781179 = 2^15 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 1^2) * 2^(-2*15) )   n = 15   d_n = 0+1i 
assign u[4'b0100] [15] = 21'h 000000;  // +0.0000152587890616 = 2^16 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 1^2) * 2^(-2*16) )   n = 16   d_n = 0+1i 
assign u[4'b0100] [16] = 21'h 000000;  // +0.0000076293945311 = 2^17 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 1^2) * 2^(-2*17) )   n = 17   d_n = 0+1i 
assign u[4'b0100] [17] = 21'h 000000;  // +0.0000038146972656 = 2^18 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 1^2) * 2^(-2*18) )   n = 18   d_n = 0+1i 
assign u[4'b0100] [18] = 21'h 000000;  // +0.0000019073486328 = 2^19 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 1^2) * 2^(-2*19) )   n = 19   d_n = 0+1i 
assign u[4'b0100] [19] = 21'h 000000;  // +0.0000009536743164 = 2^20 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 1^2) * 2^(-2*20) )   n = 20   d_n = 0+1i 
assign u[4'b0100] [20] = 21'h 000000;  // +0.0000004768371582 = 2^21 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 1^2) * 2^(-2*21) )   n = 21   d_n = 0+1i 
assign u[4'b0100] [21] = 21'h 000000;  // +0.0000002384185791 = 2^22 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 1^2) * 2^(-2*22) )   n = 22   d_n = 0+1i 
assign u[4'b0100] [22] = 21'h 000000;  // +0.0000001192092896 = 2^23 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 1^2) * 2^(-2*23) )   n = 23   d_n = 0+1i 
assign u[4'b0100] [23] = 21'h 000000;  // +0.0000000596046448 = 2^24 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 1^2) * 2^(-2*24) )   n = 24   d_n = 0+1i 
assign u[4'b0100] [24] = 21'h 000000;  // +0.0000000298023224 = 2^25 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 1^2) * 2^(-2*25) )   n = 25   d_n = 0+1i 
assign u[4'b0100] [25] = 21'h 000000;  // +0.0000000000000000 = 2^26 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 1^2) * 2^(-2*26) )   n = 26   d_n = 0+1i 
assign u[4'b0100] [26] = 21'h 000000;  // +0.0000000000000000 = 2^27 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 1^2) * 2^(-2*27) )   n = 27   d_n = 0+1i 
assign u[4'b0100] [27] = 21'h 000000;  // +0.0000000000000000 = 2^28 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 1^2) * 2^(-2*28) )   n = 28   d_n = 0+1i 
assign u[4'b0100] [28] = 21'h 000000;  // +0.0000000000000000 = 2^29 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 1^2) * 2^(-2*29) )   n = 29   d_n = 0+1i 
assign u[4'b0100] [29] = 21'h 000000;  // +0.0000000000000000 = 2^30 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 1^2) * 2^(-2*30) )   n = 30   d_n = 0+1i 
assign u[4'b0100] [30] = 21'h 000000;  // +0.0000000000000000 = 2^31 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 1^2) * 2^(-2*31) )   n = 31   d_n = 0+1i 
assign u[4'b0100] [31] = 21'h 000000;  // +0.0000000000000000 = 2^32 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 1^2) * 2^(-2*32) )   n = 32   d_n = 0+1i 
assign u[4'b0100] [32] = 21'h 000000;  // +0.0000000000000000 = 2^33 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 1^2) * 2^(-2*33) )   n = 33   d_n = 0+1i 
assign u[4'b0100] [33] = 21'h 000000;  // +0.0000000000000000 = 2^34 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 1^2) * 2^(-2*34) )   n = 34   d_n = 0+1i 
assign u[4'b0100] [34] = 21'h 000000;  // +0.0000000000000000 = 2^35 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 1^2) * 2^(-2*35) )   n = 35   d_n = 0+1i 
assign u[4'b0100] [35] = 21'h 000000;  // +0.0000000000000000 = 2^36 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 1^2) * 2^(-2*36) )   n = 36   d_n = 0+1i 
assign u[4'b0100] [36] = 21'h 000000;  // +0.0000000000000000 = 2^37 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 1^2) * 2^(-2*37) )   n = 37   d_n = 0+1i 
assign u[4'b0100] [37] = 21'h 000000;  // +0.0000000000000000 = 2^38 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 1^2) * 2^(-2*38) )   n = 38   d_n = 0+1i 
assign u[4'b0100] [38] = 21'h 000000;  // +0.0000000000000000 = 2^39 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 1^2) * 2^(-2*39) )   n = 39   d_n = 0+1i 
assign u[4'b0100] [39] = 21'h 000000;  // +0.0000000000000000 = 2^40 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 1^2) * 2^(-2*40) )   n = 40   d_n = 0+1i 
assign u[4'b0100] [40] = 21'h 000000;  // +0.0000000000000000 = 2^41 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 1^2) * 2^(-2*41) )   n = 41   d_n = 0+1i 
assign u[4'b0100] [41] = 21'h 000000;  // +0.0000000000000000 = 2^42 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 1^2) * 2^(-2*42) )   n = 42   d_n = 0+1i 
assign u[4'b0100] [42] = 21'h 000000;  // +0.0000000000000000 = 2^43 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 1^2) * 2^(-2*43) )   n = 43   d_n = 0+1i 
assign u[4'b0100] [43] = 21'h 000000;  // +0.0000000000000000 = 2^44 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 1^2) * 2^(-2*44) )   n = 44   d_n = 0+1i 
assign u[4'b0100] [44] = 21'h 000000;  // +0.0000000000000000 = 2^45 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 1^2) * 2^(-2*45) )   n = 45   d_n = 0+1i 
assign u[4'b0100] [45] = 21'h 000000;  // +0.0000000000000000 = 2^46 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 1^2) * 2^(-2*46) )   n = 46   d_n = 0+1i 
assign u[4'b0100] [46] = 21'h 000000;  // +0.0000000000000000 = 2^47 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 1^2) * 2^(-2*47) )   n = 47   d_n = 0+1i 
assign u[4'b0100] [47] = 21'h 000000;  // +0.0000000000000000 = 2^48 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 1^2) * 2^(-2*48) )   n = 48   d_n = 0+1i 
assign u[4'b0100] [48] = 21'h 000000;  // +0.0000000000000000 = 2^49 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 1^2) * 2^(-2*49) )   n = 49   d_n = 0+1i 
assign u[4'b0100] [49] = 21'h 000000;  // +0.0000000000000000 = 2^50 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 1^2) * 2^(-2*50) )   n = 50   d_n = 0+1i 
assign u[4'b0100] [50] = 21'h 000000;  // +0.0000000000000000 = 2^51 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 1^2) * 2^(-2*51) )   n = 51   d_n = 0+1i 
assign u[4'b0100] [51] = 21'h 000000;  // +0.0000000000000000 = 2^52 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 1^2) * 2^(-2*52) )   n = 52   d_n = 0+1i 
assign u[4'b0100] [52] = 21'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 1^2) * 2^(-2*53) )   n = 53   d_n = 0+1i 
assign u[4'b0100] [53] = 21'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 1^2) * 2^(-2*54) )   n = 54   d_n = 0+1i 
assign u[4'b0100] [54] = 21'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 1^2) * 2^(-2*55) )   n = 55   d_n = 0+1i 
assign u[4'b0100] [55] = 21'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 1^2) * 2^(-2*56) )   n = 56   d_n = 0+1i 
assign u[4'b0100] [56] = 21'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 1^2) * 2^(-2*57) )   n = 57   d_n = 0+1i 
assign u[4'b0100] [57] = 21'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 1^2) * 2^(-2*58) )   n = 58   d_n = 0+1i 
assign u[4'b0100] [58] = 21'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 1^2) * 2^(-2*59) )   n = 59   d_n = 0+1i 
assign u[4'b0100] [59] = 21'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 1^2) * 2^(-2*60) )   n = 60   d_n = 0+1i 
assign u[4'b0100] [60] = 21'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 1^2) * 2^(-2*61) )   n = 61   d_n = 0+1i 
assign u[4'b0100] [61] = 21'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 1^2) * 2^(-2*62) )   n = 62   d_n = 0+1i 
assign u[4'b0100] [62] = 21'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 1^2) * 2^(-2*63) )   n = 63   d_n = 0+1i 
assign u[4'b0100] [63] = 21'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 1^2) * 2^(-2*64) )   n = 64   d_n = 0+1i 
assign u[4'b0101] [00] = 21'h 000754;  // +1.8325814637483104 = 2^ 1 * ln( 1 +  1 * 2^(- 1+1) + ( 1^2+ 1^2) * 2^(-2* 1) )   n =  1   d_n = 1+1i 
assign u[4'b0101] [01] = 21'h 0007C4;  // +1.9420312631268026 = 2^ 2 * ln( 1 +  1 * 2^(- 2+1) + ( 1^2+ 1^2) * 2^(-2* 2) )   n =  2   d_n = 1+1i 
assign u[4'b0101] [02] = 21'h 0007EE;  // +1.9826893112366513 = 2^ 3 * ln( 1 +  1 * 2^(- 3+1) + ( 1^2+ 1^2) * 2^(-2* 3) )   n =  3   d_n = 1+1i 
assign u[4'b0101] [03] = 21'h 0007FB;  // +1.9952556560153185 = 2^ 4 * ln( 1 +  1 * 2^(- 4+1) + ( 1^2+ 1^2) * 2^(-2* 4) )   n =  4   d_n = 1+1i 
assign u[4'b0101] [04] = 21'h 0007FE;  // +1.9987574279595595 = 2^ 5 * ln( 1 +  1 * 2^(- 5+1) + ( 1^2+ 1^2) * 2^(-2* 5) )   n =  5   d_n = 1+1i 
assign u[4'b0101] [05] = 21'h 0007FF;  // +1.9996820132261188 = 2^ 6 * ln( 1 +  1 * 2^(- 6+1) + ( 1^2+ 1^2) * 2^(-2* 6) )   n =  6   d_n = 1+1i 
assign u[4'b0101] [06] = 21'h 0007FF;  // +1.9999195675060046 = 2^ 7 * ln( 1 +  1 * 2^(- 7+1) + ( 1^2+ 1^2) * 2^(-2* 7) )   n =  7   d_n = 1+1i 
assign u[4'b0101] [07] = 21'h 0007FF;  // +1.9999797737846823 = 2^ 8 * ln( 1 +  1 * 2^(- 8+1) + ( 1^2+ 1^2) * 2^(-2* 8) )   n =  8   d_n = 1+1i 
assign u[4'b0101] [08] = 21'h 0007FF;  // +1.9999949286148679 = 2^ 9 * ln( 1 +  1 * 2^(- 9+1) + ( 1^2+ 1^2) * 2^(-2* 9) )   n =  9   d_n = 1+1i 
assign u[4'b0101] [09] = 21'h 0007FF;  // +1.9999987302952080 = 2^10 * ln( 1 +  1 * 2^(-10+1) + ( 1^2+ 1^2) * 2^(-2*10) )   n = 10   d_n = 1+1i 
assign u[4'b0101] [10] = 21'h 0007FF;  // +1.9999996823413151 = 2^11 * ln( 1 +  1 * 2^(-11+1) + ( 1^2+ 1^2) * 2^(-2*11) )   n = 11   d_n = 1+1i 
assign u[4'b0101] [11] = 21'h 0007FF;  // +1.9999999205562393 = 2^12 * ln( 1 +  1 * 2^(-12+1) + ( 1^2+ 1^2) * 2^(-2*12) )   n = 12   d_n = 1+1i 
assign u[4'b0101] [12] = 21'h 0007FF;  // +1.9999999801340587 = 2^13 * ln( 1 +  1 * 2^(-13+1) + ( 1^2+ 1^2) * 2^(-2*13) )   n = 13   d_n = 1+1i 
assign u[4'b0101] [13] = 21'h 0007FF;  // +1.9999999950332306 = 2^14 * ln( 1 +  1 * 2^(-14+1) + ( 1^2+ 1^2) * 2^(-2*14) )   n = 14   d_n = 1+1i 
assign u[4'b0101] [14] = 21'h 0007FF;  // +1.9999999987582722 = 2^15 * ln( 1 +  1 * 2^(-15+1) + ( 1^2+ 1^2) * 2^(-2*15) )   n = 15   d_n = 1+1i 
assign u[4'b0101] [15] = 21'h 0007FF;  // +1.9999999996895637 = 2^16 * ln( 1 +  1 * 2^(-16+1) + ( 1^2+ 1^2) * 2^(-2*16) )   n = 16   d_n = 1+1i 
assign u[4'b0101] [16] = 21'h 0007FF;  // +1.9999999999223903 = 2^17 * ln( 1 +  1 * 2^(-17+1) + ( 1^2+ 1^2) * 2^(-2*17) )   n = 17   d_n = 1+1i 
assign u[4'b0101] [17] = 21'h 0007FF;  // +1.9999999999951494 = 2^18 * ln( 1 +  1 * 2^(-18+1) + ( 1^2+ 1^2) * 2^(-2*18) )   n = 18   d_n = 1+1i 
assign u[4'b0101] [18] = 21'h 0007FF;  // +1.9999999999987874 = 2^19 * ln( 1 +  1 * 2^(-19+1) + ( 1^2+ 1^2) * 2^(-2*19) )   n = 19   d_n = 1+1i 
assign u[4'b0101] [19] = 21'h 0007FF;  // +1.9999999999996969 = 2^20 * ln( 1 +  1 * 2^(-20+1) + ( 1^2+ 1^2) * 2^(-2*20) )   n = 20   d_n = 1+1i 
assign u[4'b0101] [20] = 21'h 0007FF;  // +1.9999999999999243 = 2^21 * ln( 1 +  1 * 2^(-21+1) + ( 1^2+ 1^2) * 2^(-2*21) )   n = 21   d_n = 1+1i 
assign u[4'b0101] [21] = 21'h 0007FF;  // +1.9999999999999811 = 2^22 * ln( 1 +  1 * 2^(-22+1) + ( 1^2+ 1^2) * 2^(-2*22) )   n = 22   d_n = 1+1i 
assign u[4'b0101] [22] = 21'h 0007FF;  // +1.9999999999999953 = 2^23 * ln( 1 +  1 * 2^(-23+1) + ( 1^2+ 1^2) * 2^(-2*23) )   n = 23   d_n = 1+1i 
assign u[4'b0101] [23] = 21'h 0007FF;  // +1.9999999999999989 = 2^24 * ln( 1 +  1 * 2^(-24+1) + ( 1^2+ 1^2) * 2^(-2*24) )   n = 24   d_n = 1+1i 
assign u[4'b0101] [24] = 21'h 0007FF;  // +1.9999999999999998 = 2^25 * ln( 1 +  1 * 2^(-25+1) + ( 1^2+ 1^2) * 2^(-2*25) )   n = 25   d_n = 1+1i 
assign u[4'b0101] [25] = 21'h 0007FF;  // +1.9999999850988390 = 2^26 * ln( 1 +  1 * 2^(-26+1) + ( 1^2+ 1^2) * 2^(-2*26) )   n = 26   d_n = 1+1i 
assign u[4'b0101] [26] = 21'h 0007FF;  // +1.9999999925494194 = 2^27 * ln( 1 +  1 * 2^(-27+1) + ( 1^2+ 1^2) * 2^(-2*27) )   n = 27   d_n = 1+1i 
assign u[4'b0101] [27] = 21'h 0007FF;  // +1.9999999962747097 = 2^28 * ln( 1 +  1 * 2^(-28+1) + ( 1^2+ 1^2) * 2^(-2*28) )   n = 28   d_n = 1+1i 
assign u[4'b0101] [28] = 21'h 0007FF;  // +1.9999999981373549 = 2^29 * ln( 1 +  1 * 2^(-29+1) + ( 1^2+ 1^2) * 2^(-2*29) )   n = 29   d_n = 1+1i 
assign u[4'b0101] [29] = 21'h 0007FF;  // +1.9999999990686774 = 2^30 * ln( 1 +  1 * 2^(-30+1) + ( 1^2+ 1^2) * 2^(-2*30) )   n = 30   d_n = 1+1i 
assign u[4'b0101] [30] = 21'h 0007FF;  // +1.9999999995343387 = 2^31 * ln( 1 +  1 * 2^(-31+1) + ( 1^2+ 1^2) * 2^(-2*31) )   n = 31   d_n = 1+1i 
assign u[4'b0101] [31] = 21'h 0007FF;  // +1.9999999997671694 = 2^32 * ln( 1 +  1 * 2^(-32+1) + ( 1^2+ 1^2) * 2^(-2*32) )   n = 32   d_n = 1+1i 
assign u[4'b0101] [32] = 21'h 0007FF;  // +1.9999999998835847 = 2^33 * ln( 1 +  1 * 2^(-33+1) + ( 1^2+ 1^2) * 2^(-2*33) )   n = 33   d_n = 1+1i 
assign u[4'b0101] [33] = 21'h 0007FF;  // +1.9999999999417923 = 2^34 * ln( 1 +  1 * 2^(-34+1) + ( 1^2+ 1^2) * 2^(-2*34) )   n = 34   d_n = 1+1i 
assign u[4'b0101] [34] = 21'h 0007FF;  // +1.9999999999708962 = 2^35 * ln( 1 +  1 * 2^(-35+1) + ( 1^2+ 1^2) * 2^(-2*35) )   n = 35   d_n = 1+1i 
assign u[4'b0101] [35] = 21'h 0007FF;  // +1.9999999999854481 = 2^36 * ln( 1 +  1 * 2^(-36+1) + ( 1^2+ 1^2) * 2^(-2*36) )   n = 36   d_n = 1+1i 
assign u[4'b0101] [36] = 21'h 0007FF;  // +1.9999999999927240 = 2^37 * ln( 1 +  1 * 2^(-37+1) + ( 1^2+ 1^2) * 2^(-2*37) )   n = 37   d_n = 1+1i 
assign u[4'b0101] [37] = 21'h 0007FF;  // +1.9999999999963620 = 2^38 * ln( 1 +  1 * 2^(-38+1) + ( 1^2+ 1^2) * 2^(-2*38) )   n = 38   d_n = 1+1i 
assign u[4'b0101] [38] = 21'h 0007FF;  // +1.9999999999981810 = 2^39 * ln( 1 +  1 * 2^(-39+1) + ( 1^2+ 1^2) * 2^(-2*39) )   n = 39   d_n = 1+1i 
assign u[4'b0101] [39] = 21'h 0007FF;  // +1.9999999999990905 = 2^40 * ln( 1 +  1 * 2^(-40+1) + ( 1^2+ 1^2) * 2^(-2*40) )   n = 40   d_n = 1+1i 
assign u[4'b0101] [40] = 21'h 0007FF;  // +1.9999999999995453 = 2^41 * ln( 1 +  1 * 2^(-41+1) + ( 1^2+ 1^2) * 2^(-2*41) )   n = 41   d_n = 1+1i 
assign u[4'b0101] [41] = 21'h 0007FF;  // +1.9999999999997726 = 2^42 * ln( 1 +  1 * 2^(-42+1) + ( 1^2+ 1^2) * 2^(-2*42) )   n = 42   d_n = 1+1i 
assign u[4'b0101] [42] = 21'h 0007FF;  // +1.9999999999998863 = 2^43 * ln( 1 +  1 * 2^(-43+1) + ( 1^2+ 1^2) * 2^(-2*43) )   n = 43   d_n = 1+1i 
assign u[4'b0101] [43] = 21'h 0007FF;  // +1.9999999999999432 = 2^44 * ln( 1 +  1 * 2^(-44+1) + ( 1^2+ 1^2) * 2^(-2*44) )   n = 44   d_n = 1+1i 
assign u[4'b0101] [44] = 21'h 0007FF;  // +1.9999999999999716 = 2^45 * ln( 1 +  1 * 2^(-45+1) + ( 1^2+ 1^2) * 2^(-2*45) )   n = 45   d_n = 1+1i 
assign u[4'b0101] [45] = 21'h 0007FF;  // +1.9999999999999858 = 2^46 * ln( 1 +  1 * 2^(-46+1) + ( 1^2+ 1^2) * 2^(-2*46) )   n = 46   d_n = 1+1i 
assign u[4'b0101] [46] = 21'h 0007FF;  // +1.9999999999999929 = 2^47 * ln( 1 +  1 * 2^(-47+1) + ( 1^2+ 1^2) * 2^(-2*47) )   n = 47   d_n = 1+1i 
assign u[4'b0101] [47] = 21'h 0007FF;  // +1.9999999999999964 = 2^48 * ln( 1 +  1 * 2^(-48+1) + ( 1^2+ 1^2) * 2^(-2*48) )   n = 48   d_n = 1+1i 
assign u[4'b0101] [48] = 21'h 0007FF;  // +1.9999999999999982 = 2^49 * ln( 1 +  1 * 2^(-49+1) + ( 1^2+ 1^2) * 2^(-2*49) )   n = 49   d_n = 1+1i 
assign u[4'b0101] [49] = 21'h 0007FF;  // +1.9999999999999991 = 2^50 * ln( 1 +  1 * 2^(-50+1) + ( 1^2+ 1^2) * 2^(-2*50) )   n = 50   d_n = 1+1i 
assign u[4'b0101] [50] = 21'h 0007FF;  // +1.9999999999999996 = 2^51 * ln( 1 +  1 * 2^(-51+1) + ( 1^2+ 1^2) * 2^(-2*51) )   n = 51   d_n = 1+1i 
assign u[4'b0101] [51] = 21'h 0007FF;  // +1.9999999999999998 = 2^52 * ln( 1 +  1 * 2^(-52+1) + ( 1^2+ 1^2) * 2^(-2*52) )   n = 52   d_n = 1+1i 
assign u[4'b0101] [52] = 21'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  1 * 2^(-53+1) + ( 1^2+ 1^2) * 2^(-2*53) )   n = 53   d_n = 1+1i 
assign u[4'b0101] [53] = 21'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  1 * 2^(-54+1) + ( 1^2+ 1^2) * 2^(-2*54) )   n = 54   d_n = 1+1i 
assign u[4'b0101] [54] = 21'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  1 * 2^(-55+1) + ( 1^2+ 1^2) * 2^(-2*55) )   n = 55   d_n = 1+1i 
assign u[4'b0101] [55] = 21'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  1 * 2^(-56+1) + ( 1^2+ 1^2) * 2^(-2*56) )   n = 56   d_n = 1+1i 
assign u[4'b0101] [56] = 21'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  1 * 2^(-57+1) + ( 1^2+ 1^2) * 2^(-2*57) )   n = 57   d_n = 1+1i 
assign u[4'b0101] [57] = 21'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  1 * 2^(-58+1) + ( 1^2+ 1^2) * 2^(-2*58) )   n = 58   d_n = 1+1i 
assign u[4'b0101] [58] = 21'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  1 * 2^(-59+1) + ( 1^2+ 1^2) * 2^(-2*59) )   n = 59   d_n = 1+1i 
assign u[4'b0101] [59] = 21'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  1 * 2^(-60+1) + ( 1^2+ 1^2) * 2^(-2*60) )   n = 60   d_n = 1+1i 
assign u[4'b0101] [60] = 21'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  1 * 2^(-61+1) + ( 1^2+ 1^2) * 2^(-2*61) )   n = 61   d_n = 1+1i 
assign u[4'b0101] [61] = 21'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  1 * 2^(-62+1) + ( 1^2+ 1^2) * 2^(-2*62) )   n = 62   d_n = 1+1i 
assign u[4'b0101] [62] = 21'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  1 * 2^(-63+1) + ( 1^2+ 1^2) * 2^(-2*63) )   n = 63   d_n = 1+1i 
assign u[4'b0101] [63] = 21'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  1 * 2^(-64+1) + ( 1^2+ 1^2) * 2^(-2*64) )   n = 64   d_n = 1+1i 
assign u[4'b0110] [00] = 21'h 0001C8;  // +0.4462871026284197 = 2^ 1 * ln( 1 +  0 * 2^(- 1+1) + ( 0^2+ 1^2) * 2^(-2* 1) )   n =  1   d_n = 0+1i 
assign u[4'b0110] [01] = 21'h 0000F8;  // +0.2424984872657394 = 2^ 2 * ln( 1 +  0 * 2^(- 2+1) + ( 0^2+ 1^2) * 2^(-2* 2) )   n =  2   d_n = 0+1i 
assign u[4'b0110] [02] = 21'h 00007F;  // +0.1240334922877210 = 2^ 3 * ln( 1 +  0 * 2^(- 3+1) + ( 0^2+ 1^2) * 2^(-2* 3) )   n =  3   d_n = 0+1i 
assign u[4'b0110] [03] = 21'h 00003F;  // +0.0623782466505195 = 2^ 4 * ln( 1 +  0 * 2^(- 4+1) + ( 0^2+ 1^2) * 2^(-2* 4) )   n =  4   d_n = 0+1i 
assign u[4'b0110] [04] = 21'h 00001F;  // +0.0312347511377731 = 2^ 5 * ln( 1 +  0 * 2^(- 5+1) + ( 0^2+ 1^2) * 2^(-2* 5) )   n =  5   d_n = 0+1i 
assign u[4'b0110] [05] = 21'h 00000F;  // +0.0156230929617406 = 2^ 6 * ln( 1 +  0 * 2^(- 6+1) + ( 0^2+ 1^2) * 2^(-2* 6) )   n =  6   d_n = 0+1i 
assign u[4'b0110] [06] = 21'h 000007;  // +0.0078122615911219 = 2^ 7 * ln( 1 +  0 * 2^(- 7+1) + ( 0^2+ 1^2) * 2^(-2* 7) )   n =  7   d_n = 0+1i 
assign u[4'b0110] [07] = 21'h 000003;  // +0.0039062201979808 = 2^ 8 * ln( 1 +  0 * 2^(- 8+1) + ( 0^2+ 1^2) * 2^(-2* 8) )   n =  8   d_n = 0+1i 
assign u[4'b0110] [08] = 21'h 000001;  // +0.0019531212747156 = 2^ 9 * ln( 1 +  0 * 2^(- 9+1) + ( 0^2+ 1^2) * 2^(-2* 9) )   n =  9   d_n = 0+1i 
assign u[4'b0110] [09] = 21'h 000000;  // +0.0009765620343389 = 2^10 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 1^2) * 2^(-2*10) )   n = 10   d_n = 0+1i 
assign u[4'b0110] [10] = 21'h 000000;  // +0.0004882811917923 = 2^11 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 1^2) * 2^(-2*11) )   n = 11   d_n = 0+1i 
assign u[4'b0110] [11] = 21'h 000000;  // +0.0002441406177240 = 2^12 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 1^2) * 2^(-2*12) )   n = 12   d_n = 0+1i 
assign u[4'b0110] [12] = 21'h 000000;  // +0.0001220703120453 = 2^13 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 1^2) * 2^(-2*13) )   n = 13   d_n = 0+1i 
assign u[4'b0110] [13] = 21'h 000000;  // +0.0000610351561932 = 2^14 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 1^2) * 2^(-2*14) )   n = 14   d_n = 0+1i 
assign u[4'b0110] [14] = 21'h 000000;  // +0.0000305175781179 = 2^15 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 1^2) * 2^(-2*15) )   n = 15   d_n = 0+1i 
assign u[4'b0110] [15] = 21'h 000000;  // +0.0000152587890616 = 2^16 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 1^2) * 2^(-2*16) )   n = 16   d_n = 0+1i 
assign u[4'b0110] [16] = 21'h 000000;  // +0.0000076293945311 = 2^17 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 1^2) * 2^(-2*17) )   n = 17   d_n = 0+1i 
assign u[4'b0110] [17] = 21'h 000000;  // +0.0000038146972656 = 2^18 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 1^2) * 2^(-2*18) )   n = 18   d_n = 0+1i 
assign u[4'b0110] [18] = 21'h 000000;  // +0.0000019073486328 = 2^19 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 1^2) * 2^(-2*19) )   n = 19   d_n = 0+1i 
assign u[4'b0110] [19] = 21'h 000000;  // +0.0000009536743164 = 2^20 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 1^2) * 2^(-2*20) )   n = 20   d_n = 0+1i 
assign u[4'b0110] [20] = 21'h 000000;  // +0.0000004768371582 = 2^21 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 1^2) * 2^(-2*21) )   n = 21   d_n = 0+1i 
assign u[4'b0110] [21] = 21'h 000000;  // +0.0000002384185791 = 2^22 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 1^2) * 2^(-2*22) )   n = 22   d_n = 0+1i 
assign u[4'b0110] [22] = 21'h 000000;  // +0.0000001192092896 = 2^23 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 1^2) * 2^(-2*23) )   n = 23   d_n = 0+1i 
assign u[4'b0110] [23] = 21'h 000000;  // +0.0000000596046448 = 2^24 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 1^2) * 2^(-2*24) )   n = 24   d_n = 0+1i 
assign u[4'b0110] [24] = 21'h 000000;  // +0.0000000298023224 = 2^25 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 1^2) * 2^(-2*25) )   n = 25   d_n = 0+1i 
assign u[4'b0110] [25] = 21'h 000000;  // +0.0000000000000000 = 2^26 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 1^2) * 2^(-2*26) )   n = 26   d_n = 0+1i 
assign u[4'b0110] [26] = 21'h 000000;  // +0.0000000000000000 = 2^27 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 1^2) * 2^(-2*27) )   n = 27   d_n = 0+1i 
assign u[4'b0110] [27] = 21'h 000000;  // +0.0000000000000000 = 2^28 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 1^2) * 2^(-2*28) )   n = 28   d_n = 0+1i 
assign u[4'b0110] [28] = 21'h 000000;  // +0.0000000000000000 = 2^29 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 1^2) * 2^(-2*29) )   n = 29   d_n = 0+1i 
assign u[4'b0110] [29] = 21'h 000000;  // +0.0000000000000000 = 2^30 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 1^2) * 2^(-2*30) )   n = 30   d_n = 0+1i 
assign u[4'b0110] [30] = 21'h 000000;  // +0.0000000000000000 = 2^31 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 1^2) * 2^(-2*31) )   n = 31   d_n = 0+1i 
assign u[4'b0110] [31] = 21'h 000000;  // +0.0000000000000000 = 2^32 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 1^2) * 2^(-2*32) )   n = 32   d_n = 0+1i 
assign u[4'b0110] [32] = 21'h 000000;  // +0.0000000000000000 = 2^33 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 1^2) * 2^(-2*33) )   n = 33   d_n = 0+1i 
assign u[4'b0110] [33] = 21'h 000000;  // +0.0000000000000000 = 2^34 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 1^2) * 2^(-2*34) )   n = 34   d_n = 0+1i 
assign u[4'b0110] [34] = 21'h 000000;  // +0.0000000000000000 = 2^35 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 1^2) * 2^(-2*35) )   n = 35   d_n = 0+1i 
assign u[4'b0110] [35] = 21'h 000000;  // +0.0000000000000000 = 2^36 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 1^2) * 2^(-2*36) )   n = 36   d_n = 0+1i 
assign u[4'b0110] [36] = 21'h 000000;  // +0.0000000000000000 = 2^37 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 1^2) * 2^(-2*37) )   n = 37   d_n = 0+1i 
assign u[4'b0110] [37] = 21'h 000000;  // +0.0000000000000000 = 2^38 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 1^2) * 2^(-2*38) )   n = 38   d_n = 0+1i 
assign u[4'b0110] [38] = 21'h 000000;  // +0.0000000000000000 = 2^39 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 1^2) * 2^(-2*39) )   n = 39   d_n = 0+1i 
assign u[4'b0110] [39] = 21'h 000000;  // +0.0000000000000000 = 2^40 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 1^2) * 2^(-2*40) )   n = 40   d_n = 0+1i 
assign u[4'b0110] [40] = 21'h 000000;  // +0.0000000000000000 = 2^41 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 1^2) * 2^(-2*41) )   n = 41   d_n = 0+1i 
assign u[4'b0110] [41] = 21'h 000000;  // +0.0000000000000000 = 2^42 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 1^2) * 2^(-2*42) )   n = 42   d_n = 0+1i 
assign u[4'b0110] [42] = 21'h 000000;  // +0.0000000000000000 = 2^43 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 1^2) * 2^(-2*43) )   n = 43   d_n = 0+1i 
assign u[4'b0110] [43] = 21'h 000000;  // +0.0000000000000000 = 2^44 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 1^2) * 2^(-2*44) )   n = 44   d_n = 0+1i 
assign u[4'b0110] [44] = 21'h 000000;  // +0.0000000000000000 = 2^45 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 1^2) * 2^(-2*45) )   n = 45   d_n = 0+1i 
assign u[4'b0110] [45] = 21'h 000000;  // +0.0000000000000000 = 2^46 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 1^2) * 2^(-2*46) )   n = 46   d_n = 0+1i 
assign u[4'b0110] [46] = 21'h 000000;  // +0.0000000000000000 = 2^47 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 1^2) * 2^(-2*47) )   n = 47   d_n = 0+1i 
assign u[4'b0110] [47] = 21'h 000000;  // +0.0000000000000000 = 2^48 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 1^2) * 2^(-2*48) )   n = 48   d_n = 0+1i 
assign u[4'b0110] [48] = 21'h 000000;  // +0.0000000000000000 = 2^49 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 1^2) * 2^(-2*49) )   n = 49   d_n = 0+1i 
assign u[4'b0110] [49] = 21'h 000000;  // +0.0000000000000000 = 2^50 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 1^2) * 2^(-2*50) )   n = 50   d_n = 0+1i 
assign u[4'b0110] [50] = 21'h 000000;  // +0.0000000000000000 = 2^51 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 1^2) * 2^(-2*51) )   n = 51   d_n = 0+1i 
assign u[4'b0110] [51] = 21'h 000000;  // +0.0000000000000000 = 2^52 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 1^2) * 2^(-2*52) )   n = 52   d_n = 0+1i 
assign u[4'b0110] [52] = 21'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 1^2) * 2^(-2*53) )   n = 53   d_n = 0+1i 
assign u[4'b0110] [53] = 21'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 1^2) * 2^(-2*54) )   n = 54   d_n = 0+1i 
assign u[4'b0110] [54] = 21'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 1^2) * 2^(-2*55) )   n = 55   d_n = 0+1i 
assign u[4'b0110] [55] = 21'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 1^2) * 2^(-2*56) )   n = 56   d_n = 0+1i 
assign u[4'b0110] [56] = 21'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 1^2) * 2^(-2*57) )   n = 57   d_n = 0+1i 
assign u[4'b0110] [57] = 21'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 1^2) * 2^(-2*58) )   n = 58   d_n = 0+1i 
assign u[4'b0110] [58] = 21'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 1^2) * 2^(-2*59) )   n = 59   d_n = 0+1i 
assign u[4'b0110] [59] = 21'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 1^2) * 2^(-2*60) )   n = 60   d_n = 0+1i 
assign u[4'b0110] [60] = 21'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 1^2) * 2^(-2*61) )   n = 61   d_n = 0+1i 
assign u[4'b0110] [61] = 21'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 1^2) * 2^(-2*62) )   n = 62   d_n = 0+1i 
assign u[4'b0110] [62] = 21'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 1^2) * 2^(-2*63) )   n = 63   d_n = 0+1i 
assign u[4'b0110] [63] = 21'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 1^2) * 2^(-2*64) )   n = 64   d_n = 0+1i 
assign u[4'b0111] [00] = 21'h 1FFA74;  // -1.3862943611198904 = 2^ 1 * ln( 1 + -1 * 2^(- 1+1) + (-1^2+ 1^2) * 2^(-2* 1) )   n =  1   d_n = -1+1i 
assign u[4'b0111] [01] = 21'h 1FF87A;  // -1.8800145169829416 = 2^ 2 * ln( 1 + -1 * 2^(- 2+1) + (-1^2+ 1^2) * 2^(-2* 2) )   n =  2   d_n = -1+1i 
assign u[4'b0111] [02] = 21'h 1FF819;  // -1.9748806234522058 = 2^ 3 * ln( 1 + -1 * 2^(- 3+1) + (-1^2+ 1^2) * 2^(-2* 3) )   n =  3   d_n = -1+1i 
assign u[4'b0111] [03] = 21'h 1FF805;  // -1.9942791233164259 = 2^ 4 * ln( 1 + -1 * 2^(- 4+1) + (-1^2+ 1^2) * 2^(-2* 4) )   n =  4   d_n = -1+1i 
assign u[4'b0111] [04] = 21'h 1FF801;  // -1.9986353578798890 = 2^ 5 * ln( 1 + -1 * 2^(- 5+1) + (-1^2+ 1^2) * 2^(-2* 5) )   n =  5   d_n = -1+1i 
assign u[4'b0111] [05] = 21'h 1FF800;  // -1.9996667544388824 = 2^ 6 * ln( 1 + -1 * 2^(- 6+1) + (-1^2+ 1^2) * 2^(-2* 6) )   n =  6   d_n = -1+1i 
assign u[4'b0111] [06] = 21'h 1FF800;  // -1.9999176601574109 = 2^ 7 * ln( 1 + -1 * 2^(- 7+1) + (-1^2+ 1^2) * 2^(-2* 7) )   n =  7   d_n = -1+1i 
assign u[4'b0111] [07] = 21'h 1FF800;  // -1.9999795353661032 = 2^ 8 * ln( 1 + -1 * 2^(- 8+1) + (-1^2+ 1^2) * 2^(-2* 8) )   n =  8   d_n = -1+1i 
assign u[4'b0111] [08] = 21'h 1FF800;  // -1.9999948988125242 = 2^ 9 * ln( 1 + -1 * 2^(- 9+1) + (-1^2+ 1^2) * 2^(-2* 9) )   n =  9   d_n = -1+1i 
assign u[4'b0111] [09] = 21'h 1FF800;  // -1.9999987265701442 = 2^10 * ln( 1 + -1 * 2^(-10+1) + (-1^2+ 1^2) * 2^(-2*10) )   n = 10   d_n = -1+1i 
assign u[4'b0111] [10] = 21'h 1FF800;  // -1.9999996818756538 = 2^11 * ln( 1 + -1 * 2^(-11+1) + (-1^2+ 1^2) * 2^(-2*11) )   n = 11   d_n = -1+1i 
assign u[4'b0111] [11] = 21'h 1FF800;  // -1.9999999204980317 = 2^12 * ln( 1 + -1 * 2^(-12+1) + (-1^2+ 1^2) * 2^(-2*12) )   n = 12   d_n = -1+1i 
assign u[4'b0111] [12] = 21'h 1FF800;  // -1.9999999801276920 = 2^13 * ln( 1 + -1 * 2^(-13+1) + (-1^2+ 1^2) * 2^(-2*13) )   n = 13   d_n = -1+1i 
assign u[4'b0111] [13] = 21'h 1FF800;  // -1.9999999950326621 = 2^14 * ln( 1 + -1 * 2^(-14+1) + (-1^2+ 1^2) * 2^(-2*14) )   n = 14   d_n = -1+1i 
assign u[4'b0111] [14] = 21'h 1FF800;  // -1.9999999987582011 = 2^15 * ln( 1 + -1 * 2^(-15+1) + (-1^2+ 1^2) * 2^(-2*15) )   n = 15   d_n = -1+1i 
assign u[4'b0111] [15] = 21'h 1FF800;  // -1.9999999996895548 = 2^16 * ln( 1 + -1 * 2^(-16+1) + (-1^2+ 1^2) * 2^(-2*16) )   n = 16   d_n = -1+1i 
assign u[4'b0111] [16] = 21'h 1FF800;  // -1.9999999999223892 = 2^17 * ln( 1 + -1 * 2^(-17+1) + (-1^2+ 1^2) * 2^(-2*17) )   n = 17   d_n = -1+1i 
assign u[4'b0111] [17] = 21'h 1FF800;  // -1.9999999999951494 = 2^18 * ln( 1 + -1 * 2^(-18+1) + (-1^2+ 1^2) * 2^(-2*18) )   n = 18   d_n = -1+1i 
assign u[4'b0111] [18] = 21'h 1FF800;  // -1.9999999999987874 = 2^19 * ln( 1 + -1 * 2^(-19+1) + (-1^2+ 1^2) * 2^(-2*19) )   n = 19   d_n = -1+1i 
assign u[4'b0111] [19] = 21'h 1FF800;  // -1.9999999999996969 = 2^20 * ln( 1 + -1 * 2^(-20+1) + (-1^2+ 1^2) * 2^(-2*20) )   n = 20   d_n = -1+1i 
assign u[4'b0111] [20] = 21'h 1FF800;  // -1.9999999999999243 = 2^21 * ln( 1 + -1 * 2^(-21+1) + (-1^2+ 1^2) * 2^(-2*21) )   n = 21   d_n = -1+1i 
assign u[4'b0111] [21] = 21'h 1FF800;  // -1.9999999999999811 = 2^22 * ln( 1 + -1 * 2^(-22+1) + (-1^2+ 1^2) * 2^(-2*22) )   n = 22   d_n = -1+1i 
assign u[4'b0111] [22] = 21'h 1FF800;  // -1.9999999999999953 = 2^23 * ln( 1 + -1 * 2^(-23+1) + (-1^2+ 1^2) * 2^(-2*23) )   n = 23   d_n = -1+1i 
assign u[4'b0111] [23] = 21'h 1FF800;  // -1.9999999999999989 = 2^24 * ln( 1 + -1 * 2^(-24+1) + (-1^2+ 1^2) * 2^(-2*24) )   n = 24   d_n = -1+1i 
assign u[4'b0111] [24] = 21'h 1FF800;  // -1.9999999999999998 = 2^25 * ln( 1 + -1 * 2^(-25+1) + (-1^2+ 1^2) * 2^(-2*25) )   n = 25   d_n = -1+1i 
assign u[4'b0111] [25] = 21'h 1FF800;  // -2.0000000000000000 = 2^26 * ln( 1 + -1 * 2^(-26+1) + (-1^2+ 1^2) * 2^(-2*26) )   n = 26   d_n = -1+1i 
assign u[4'b0111] [26] = 21'h 1FF7FF;  // -2.0000000074505806 = 2^27 * ln( 1 + -1 * 2^(-27+1) + (-1^2+ 1^2) * 2^(-2*27) )   n = 27   d_n = -1+1i 
assign u[4'b0111] [27] = 21'h 1FF7FF;  // -2.0000000037252903 = 2^28 * ln( 1 + -1 * 2^(-28+1) + (-1^2+ 1^2) * 2^(-2*28) )   n = 28   d_n = -1+1i 
assign u[4'b0111] [28] = 21'h 1FF7FF;  // -2.0000000018626451 = 2^29 * ln( 1 + -1 * 2^(-29+1) + (-1^2+ 1^2) * 2^(-2*29) )   n = 29   d_n = -1+1i 
assign u[4'b0111] [29] = 21'h 1FF7FF;  // -2.0000000009313226 = 2^30 * ln( 1 + -1 * 2^(-30+1) + (-1^2+ 1^2) * 2^(-2*30) )   n = 30   d_n = -1+1i 
assign u[4'b0111] [30] = 21'h 1FF7FF;  // -2.0000000004656613 = 2^31 * ln( 1 + -1 * 2^(-31+1) + (-1^2+ 1^2) * 2^(-2*31) )   n = 31   d_n = -1+1i 
assign u[4'b0111] [31] = 21'h 1FF7FF;  // -2.0000000002328306 = 2^32 * ln( 1 + -1 * 2^(-32+1) + (-1^2+ 1^2) * 2^(-2*32) )   n = 32   d_n = -1+1i 
assign u[4'b0111] [32] = 21'h 1FF7FF;  // -2.0000000001164153 = 2^33 * ln( 1 + -1 * 2^(-33+1) + (-1^2+ 1^2) * 2^(-2*33) )   n = 33   d_n = -1+1i 
assign u[4'b0111] [33] = 21'h 1FF7FF;  // -2.0000000000582077 = 2^34 * ln( 1 + -1 * 2^(-34+1) + (-1^2+ 1^2) * 2^(-2*34) )   n = 34   d_n = -1+1i 
assign u[4'b0111] [34] = 21'h 1FF7FF;  // -2.0000000000291038 = 2^35 * ln( 1 + -1 * 2^(-35+1) + (-1^2+ 1^2) * 2^(-2*35) )   n = 35   d_n = -1+1i 
assign u[4'b0111] [35] = 21'h 1FF7FF;  // -2.0000000000145519 = 2^36 * ln( 1 + -1 * 2^(-36+1) + (-1^2+ 1^2) * 2^(-2*36) )   n = 36   d_n = -1+1i 
assign u[4'b0111] [36] = 21'h 1FF7FF;  // -2.0000000000072760 = 2^37 * ln( 1 + -1 * 2^(-37+1) + (-1^2+ 1^2) * 2^(-2*37) )   n = 37   d_n = -1+1i 
assign u[4'b0111] [37] = 21'h 1FF7FF;  // -2.0000000000036380 = 2^38 * ln( 1 + -1 * 2^(-38+1) + (-1^2+ 1^2) * 2^(-2*38) )   n = 38   d_n = -1+1i 
assign u[4'b0111] [38] = 21'h 1FF7FF;  // -2.0000000000018190 = 2^39 * ln( 1 + -1 * 2^(-39+1) + (-1^2+ 1^2) * 2^(-2*39) )   n = 39   d_n = -1+1i 
assign u[4'b0111] [39] = 21'h 1FF7FF;  // -2.0000000000009095 = 2^40 * ln( 1 + -1 * 2^(-40+1) + (-1^2+ 1^2) * 2^(-2*40) )   n = 40   d_n = -1+1i 
assign u[4'b0111] [40] = 21'h 1FF7FF;  // -2.0000000000004547 = 2^41 * ln( 1 + -1 * 2^(-41+1) + (-1^2+ 1^2) * 2^(-2*41) )   n = 41   d_n = -1+1i 
assign u[4'b0111] [41] = 21'h 1FF7FF;  // -2.0000000000002274 = 2^42 * ln( 1 + -1 * 2^(-42+1) + (-1^2+ 1^2) * 2^(-2*42) )   n = 42   d_n = -1+1i 
assign u[4'b0111] [42] = 21'h 1FF800;  // -2.0000000000001137 = 2^43 * ln( 1 + -1 * 2^(-43+1) + (-1^2+ 1^2) * 2^(-2*43) )   n = 43   d_n = -1+1i 
assign u[4'b0111] [43] = 21'h 1FF800;  // -2.0000000000000568 = 2^44 * ln( 1 + -1 * 2^(-44+1) + (-1^2+ 1^2) * 2^(-2*44) )   n = 44   d_n = -1+1i 
assign u[4'b0111] [44] = 21'h 1FF800;  // -2.0000000000000284 = 2^45 * ln( 1 + -1 * 2^(-45+1) + (-1^2+ 1^2) * 2^(-2*45) )   n = 45   d_n = -1+1i 
assign u[4'b0111] [45] = 21'h 1FF800;  // -2.0000000000000142 = 2^46 * ln( 1 + -1 * 2^(-46+1) + (-1^2+ 1^2) * 2^(-2*46) )   n = 46   d_n = -1+1i 
assign u[4'b0111] [46] = 21'h 1FF800;  // -2.0000000000000071 = 2^47 * ln( 1 + -1 * 2^(-47+1) + (-1^2+ 1^2) * 2^(-2*47) )   n = 47   d_n = -1+1i 
assign u[4'b0111] [47] = 21'h 1FF800;  // -2.0000000000000036 = 2^48 * ln( 1 + -1 * 2^(-48+1) + (-1^2+ 1^2) * 2^(-2*48) )   n = 48   d_n = -1+1i 
assign u[4'b0111] [48] = 21'h 1FF800;  // -2.0000000000000018 = 2^49 * ln( 1 + -1 * 2^(-49+1) + (-1^2+ 1^2) * 2^(-2*49) )   n = 49   d_n = -1+1i 
assign u[4'b0111] [49] = 21'h 1FF800;  // -2.0000000000000009 = 2^50 * ln( 1 + -1 * 2^(-50+1) + (-1^2+ 1^2) * 2^(-2*50) )   n = 50   d_n = -1+1i 
assign u[4'b0111] [50] = 21'h 1FF800;  // -2.0000000000000004 = 2^51 * ln( 1 + -1 * 2^(-51+1) + (-1^2+ 1^2) * 2^(-2*51) )   n = 51   d_n = -1+1i 
assign u[4'b0111] [51] = 21'h 1FF800;  // -2.0000000000000004 = 2^52 * ln( 1 + -1 * 2^(-52+1) + (-1^2+ 1^2) * 2^(-2*52) )   n = 52   d_n = -1+1i 
assign u[4'b0111] [52] = 21'h 1FF800;  // -2.0000000000000000 = 2^53 * ln( 1 + -1 * 2^(-53+1) + (-1^2+ 1^2) * 2^(-2*53) )   n = 53   d_n = -1+1i 
assign u[4'b0111] [53] = 21'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 + -1 * 2^(-54+1) + (-1^2+ 1^2) * 2^(-2*54) )   n = 54   d_n = -1+1i 
assign u[4'b0111] [54] = 21'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 + -1 * 2^(-55+1) + (-1^2+ 1^2) * 2^(-2*55) )   n = 55   d_n = -1+1i 
assign u[4'b0111] [55] = 21'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 + -1 * 2^(-56+1) + (-1^2+ 1^2) * 2^(-2*56) )   n = 56   d_n = -1+1i 
assign u[4'b0111] [56] = 21'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 + -1 * 2^(-57+1) + (-1^2+ 1^2) * 2^(-2*57) )   n = 57   d_n = -1+1i 
assign u[4'b0111] [57] = 21'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 + -1 * 2^(-58+1) + (-1^2+ 1^2) * 2^(-2*58) )   n = 58   d_n = -1+1i 
assign u[4'b0111] [58] = 21'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 + -1 * 2^(-59+1) + (-1^2+ 1^2) * 2^(-2*59) )   n = 59   d_n = -1+1i 
assign u[4'b0111] [59] = 21'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 + -1 * 2^(-60+1) + (-1^2+ 1^2) * 2^(-2*60) )   n = 60   d_n = -1+1i 
assign u[4'b0111] [60] = 21'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 + -1 * 2^(-61+1) + (-1^2+ 1^2) * 2^(-2*61) )   n = 61   d_n = -1+1i 
assign u[4'b0111] [61] = 21'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 + -1 * 2^(-62+1) + (-1^2+ 1^2) * 2^(-2*62) )   n = 62   d_n = -1+1i 
assign u[4'b0111] [62] = 21'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 + -1 * 2^(-63+1) + (-1^2+ 1^2) * 2^(-2*63) )   n = 63   d_n = -1+1i 
assign u[4'b0111] [63] = 21'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 + -1 * 2^(-64+1) + (-1^2+ 1^2) * 2^(-2*64) )   n = 64   d_n = -1+1i 
assign u[4'b1000] [00] = 21'h 000000;  // +0.0000000000000000 = 2^ 1 * ln( 1 +  0 * 2^(- 1+1) + ( 0^2+ 0^2) * 2^(-2* 1) )   n =  1   d_n = 0 
assign u[4'b1000] [01] = 21'h 000000;  // +0.0000000000000000 = 2^ 2 * ln( 1 +  0 * 2^(- 2+1) + ( 0^2+ 0^2) * 2^(-2* 2) )   n =  2   d_n = 0 
assign u[4'b1000] [02] = 21'h 000000;  // +0.0000000000000000 = 2^ 3 * ln( 1 +  0 * 2^(- 3+1) + ( 0^2+ 0^2) * 2^(-2* 3) )   n =  3   d_n = 0 
assign u[4'b1000] [03] = 21'h 000000;  // +0.0000000000000000 = 2^ 4 * ln( 1 +  0 * 2^(- 4+1) + ( 0^2+ 0^2) * 2^(-2* 4) )   n =  4   d_n = 0 
assign u[4'b1000] [04] = 21'h 000000;  // +0.0000000000000000 = 2^ 5 * ln( 1 +  0 * 2^(- 5+1) + ( 0^2+ 0^2) * 2^(-2* 5) )   n =  5   d_n = 0 
assign u[4'b1000] [05] = 21'h 000000;  // +0.0000000000000000 = 2^ 6 * ln( 1 +  0 * 2^(- 6+1) + ( 0^2+ 0^2) * 2^(-2* 6) )   n =  6   d_n = 0 
assign u[4'b1000] [06] = 21'h 000000;  // +0.0000000000000000 = 2^ 7 * ln( 1 +  0 * 2^(- 7+1) + ( 0^2+ 0^2) * 2^(-2* 7) )   n =  7   d_n = 0 
assign u[4'b1000] [07] = 21'h 000000;  // +0.0000000000000000 = 2^ 8 * ln( 1 +  0 * 2^(- 8+1) + ( 0^2+ 0^2) * 2^(-2* 8) )   n =  8   d_n = 0 
assign u[4'b1000] [08] = 21'h 000000;  // +0.0000000000000000 = 2^ 9 * ln( 1 +  0 * 2^(- 9+1) + ( 0^2+ 0^2) * 2^(-2* 9) )   n =  9   d_n = 0 
assign u[4'b1000] [09] = 21'h 000000;  // +0.0000000000000000 = 2^10 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = 0 
assign u[4'b1000] [10] = 21'h 000000;  // +0.0000000000000000 = 2^11 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = 0 
assign u[4'b1000] [11] = 21'h 000000;  // +0.0000000000000000 = 2^12 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = 0 
assign u[4'b1000] [12] = 21'h 000000;  // +0.0000000000000000 = 2^13 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = 0 
assign u[4'b1000] [13] = 21'h 000000;  // +0.0000000000000000 = 2^14 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = 0 
assign u[4'b1000] [14] = 21'h 000000;  // +0.0000000000000000 = 2^15 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = 0 
assign u[4'b1000] [15] = 21'h 000000;  // +0.0000000000000000 = 2^16 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = 0 
assign u[4'b1000] [16] = 21'h 000000;  // +0.0000000000000000 = 2^17 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = 0 
assign u[4'b1000] [17] = 21'h 000000;  // +0.0000000000000000 = 2^18 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = 0 
assign u[4'b1000] [18] = 21'h 000000;  // +0.0000000000000000 = 2^19 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = 0 
assign u[4'b1000] [19] = 21'h 000000;  // +0.0000000000000000 = 2^20 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = 0 
assign u[4'b1000] [20] = 21'h 000000;  // +0.0000000000000000 = 2^21 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = 0 
assign u[4'b1000] [21] = 21'h 000000;  // +0.0000000000000000 = 2^22 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = 0 
assign u[4'b1000] [22] = 21'h 000000;  // +0.0000000000000000 = 2^23 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = 0 
assign u[4'b1000] [23] = 21'h 000000;  // +0.0000000000000000 = 2^24 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = 0 
assign u[4'b1000] [24] = 21'h 000000;  // +0.0000000000000000 = 2^25 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = 0 
assign u[4'b1000] [25] = 21'h 000000;  // +0.0000000000000000 = 2^26 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = 0 
assign u[4'b1000] [26] = 21'h 000000;  // +0.0000000000000000 = 2^27 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = 0 
assign u[4'b1000] [27] = 21'h 000000;  // +0.0000000000000000 = 2^28 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = 0 
assign u[4'b1000] [28] = 21'h 000000;  // +0.0000000000000000 = 2^29 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = 0 
assign u[4'b1000] [29] = 21'h 000000;  // +0.0000000000000000 = 2^30 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = 0 
assign u[4'b1000] [30] = 21'h 000000;  // +0.0000000000000000 = 2^31 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = 0 
assign u[4'b1000] [31] = 21'h 000000;  // +0.0000000000000000 = 2^32 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = 0 
assign u[4'b1000] [32] = 21'h 000000;  // +0.0000000000000000 = 2^33 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = 0 
assign u[4'b1000] [33] = 21'h 000000;  // +0.0000000000000000 = 2^34 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = 0 
assign u[4'b1000] [34] = 21'h 000000;  // +0.0000000000000000 = 2^35 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = 0 
assign u[4'b1000] [35] = 21'h 000000;  // +0.0000000000000000 = 2^36 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = 0 
assign u[4'b1000] [36] = 21'h 000000;  // +0.0000000000000000 = 2^37 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = 0 
assign u[4'b1000] [37] = 21'h 000000;  // +0.0000000000000000 = 2^38 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = 0 
assign u[4'b1000] [38] = 21'h 000000;  // +0.0000000000000000 = 2^39 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = 0 
assign u[4'b1000] [39] = 21'h 000000;  // +0.0000000000000000 = 2^40 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = 0 
assign u[4'b1000] [40] = 21'h 000000;  // +0.0000000000000000 = 2^41 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = 0 
assign u[4'b1000] [41] = 21'h 000000;  // +0.0000000000000000 = 2^42 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = 0 
assign u[4'b1000] [42] = 21'h 000000;  // +0.0000000000000000 = 2^43 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = 0 
assign u[4'b1000] [43] = 21'h 000000;  // +0.0000000000000000 = 2^44 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = 0 
assign u[4'b1000] [44] = 21'h 000000;  // +0.0000000000000000 = 2^45 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = 0 
assign u[4'b1000] [45] = 21'h 000000;  // +0.0000000000000000 = 2^46 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = 0 
assign u[4'b1000] [46] = 21'h 000000;  // +0.0000000000000000 = 2^47 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = 0 
assign u[4'b1000] [47] = 21'h 000000;  // +0.0000000000000000 = 2^48 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = 0 
assign u[4'b1000] [48] = 21'h 000000;  // +0.0000000000000000 = 2^49 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = 0 
assign u[4'b1000] [49] = 21'h 000000;  // +0.0000000000000000 = 2^50 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = 0 
assign u[4'b1000] [50] = 21'h 000000;  // +0.0000000000000000 = 2^51 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = 0 
assign u[4'b1000] [51] = 21'h 000000;  // +0.0000000000000000 = 2^52 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = 0 
assign u[4'b1000] [52] = 21'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = 0 
assign u[4'b1000] [53] = 21'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = 0 
assign u[4'b1000] [54] = 21'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = 0 
assign u[4'b1000] [55] = 21'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = 0 
assign u[4'b1000] [56] = 21'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = 0 
assign u[4'b1000] [57] = 21'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = 0 
assign u[4'b1000] [58] = 21'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = 0 
assign u[4'b1000] [59] = 21'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = 0 
assign u[4'b1000] [60] = 21'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = 0 
assign u[4'b1000] [61] = 21'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = 0 
assign u[4'b1000] [62] = 21'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = 0 
assign u[4'b1000] [63] = 21'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = 0 
assign u[4'b1001] [00] = 21'h 00067C;  // +1.6218604324326575 = 2^ 1 * ln( 1 +  1 * 2^(- 1+1) + ( 1^2+ 0^2) * 2^(-2* 1) )   n =  1   d_n = 1 
assign u[4'b1001] [01] = 21'h 000723;  // +1.7851484105136781 = 2^ 2 * ln( 1 +  1 * 2^(- 2+1) + ( 1^2+ 0^2) * 2^(-2* 2) )   n =  2   d_n = 1 
assign u[4'b1001] [02] = 21'h 000789;  // +1.8845285705021353 = 2^ 3 * ln( 1 +  1 * 2^(- 3+1) + ( 1^2+ 0^2) * 2^(-2* 3) )   n =  3   d_n = 1 
assign u[4'b1001] [03] = 21'h 0007C2;  // +1.9399878981259149 = 2^ 4 * ln( 1 +  1 * 2^(- 4+1) + ( 1^2+ 0^2) * 2^(-2* 4) )   n =  4   d_n = 1 
assign u[4'b1001] [04] = 21'h 0007E0;  // +1.9693861546722360 = 2^ 5 * ln( 1 +  1 * 2^(- 5+1) + ( 1^2+ 0^2) * 2^(-2* 5) )   n =  5   d_n = 1 
assign u[4'b1001] [05] = 21'h 0007F0;  // +1.9845358766035526 = 2^ 6 * ln( 1 +  1 * 2^(- 6+1) + ( 1^2+ 0^2) * 2^(-2* 6) )   n =  6   d_n = 1 
assign u[4'b1001] [06] = 21'h 0007F8;  // +1.9922279531660669 = 2^ 7 * ln( 1 +  1 * 2^(- 7+1) + ( 1^2+ 0^2) * 2^(-2* 7) )   n =  7   d_n = 1 
assign u[4'b1001] [07] = 21'h 0007FC;  // +1.9961038928165493 = 2^ 8 * ln( 1 +  1 * 2^(- 8+1) + ( 1^2+ 0^2) * 2^(-2* 8) )   n =  8   d_n = 1 
assign u[4'b1001] [08] = 21'h 0007FE;  // +1.9980494144120313 = 2^ 9 * ln( 1 +  1 * 2^(- 9+1) + ( 1^2+ 0^2) * 2^(-2* 9) )   n =  9   d_n = 1 
assign u[4'b1001] [09] = 21'h 0007FF;  // +1.9990240728175799 = 2^10 * ln( 1 +  1 * 2^(-10+1) + ( 1^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = 1 
assign u[4'b1001] [10] = 21'h 0007FF;  // +1.9995118776375345 = 2^11 * ln( 1 +  1 * 2^(-11+1) + ( 1^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = 1 
assign u[4'b1001] [11] = 21'h 0007FF;  // +1.9997558991041553 = 2^12 * ln( 1 +  1 * 2^(-12+1) + ( 1^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = 1 
assign u[4'b1001] [12] = 21'h 0007FF;  // +1.9998779396206980 = 2^13 * ln( 1 +  1 * 2^(-13+1) + ( 1^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = 1 
assign u[4'b1001] [13] = 21'h 0007FF;  // +1.9999389673271633 = 2^14 * ln( 1 +  1 * 2^(-14+1) + ( 1^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = 1 
assign u[4'b1001] [14] = 21'h 0007FF;  // +1.9999694830427426 = 2^15 * ln( 1 +  1 * 2^(-15+1) + ( 1^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = 1 
assign u[4'b1001] [15] = 21'h 0007FF;  // +1.9999847413661562 = 2^16 * ln( 1 +  1 * 2^(-16+1) + ( 1^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = 1 
assign u[4'b1001] [16] = 21'h 0007FF;  // +1.9999923706442737 = 2^17 * ln( 1 +  1 * 2^(-17+1) + ( 1^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = 1 
assign u[4'b1001] [17] = 21'h 0007FF;  // +1.9999961853124357 = 2^18 * ln( 1 +  1 * 2^(-18+1) + ( 1^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = 1 
assign u[4'b1001] [18] = 21'h 0007FF;  // +1.9999980926537926 = 2^19 * ln( 1 +  1 * 2^(-19+1) + ( 1^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = 1 
assign u[4'b1001] [19] = 21'h 0007FF;  // +1.9999990463262900 = 2^20 * ln( 1 +  1 * 2^(-20+1) + ( 1^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = 1 
assign u[4'b1001] [20] = 21'h 0007FF;  // +1.9999995231629935 = 2^21 * ln( 1 +  1 * 2^(-21+1) + ( 1^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = 1 
assign u[4'b1001] [21] = 21'h 0007FF;  // +1.9999997615814589 = 2^22 * ln( 1 +  1 * 2^(-22+1) + ( 1^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = 1 
assign u[4'b1001] [22] = 21'h 0007FF;  // +1.9999998807907200 = 2^23 * ln( 1 +  1 * 2^(-23+1) + ( 1^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = 1 
assign u[4'b1001] [23] = 21'h 0007FF;  // +1.9999999403953577 = 2^24 * ln( 1 +  1 * 2^(-24+1) + ( 1^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = 1 
assign u[4'b1001] [24] = 21'h 0007FF;  // +1.9999999701976783 = 2^25 * ln( 1 +  1 * 2^(-25+1) + ( 1^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = 1 
assign u[4'b1001] [25] = 21'h 0007FF;  // +1.9999999850988390 = 2^26 * ln( 1 +  1 * 2^(-26+1) + ( 1^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = 1 
assign u[4'b1001] [26] = 21'h 0007FF;  // +1.9999999925494194 = 2^27 * ln( 1 +  1 * 2^(-27+1) + ( 1^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = 1 
assign u[4'b1001] [27] = 21'h 0007FF;  // +1.9999999962747097 = 2^28 * ln( 1 +  1 * 2^(-28+1) + ( 1^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = 1 
assign u[4'b1001] [28] = 21'h 0007FF;  // +1.9999999981373549 = 2^29 * ln( 1 +  1 * 2^(-29+1) + ( 1^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = 1 
assign u[4'b1001] [29] = 21'h 0007FF;  // +1.9999999990686774 = 2^30 * ln( 1 +  1 * 2^(-30+1) + ( 1^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = 1 
assign u[4'b1001] [30] = 21'h 0007FF;  // +1.9999999995343387 = 2^31 * ln( 1 +  1 * 2^(-31+1) + ( 1^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = 1 
assign u[4'b1001] [31] = 21'h 0007FF;  // +1.9999999997671694 = 2^32 * ln( 1 +  1 * 2^(-32+1) + ( 1^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = 1 
assign u[4'b1001] [32] = 21'h 0007FF;  // +1.9999999998835847 = 2^33 * ln( 1 +  1 * 2^(-33+1) + ( 1^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = 1 
assign u[4'b1001] [33] = 21'h 0007FF;  // +1.9999999999417923 = 2^34 * ln( 1 +  1 * 2^(-34+1) + ( 1^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = 1 
assign u[4'b1001] [34] = 21'h 0007FF;  // +1.9999999999708962 = 2^35 * ln( 1 +  1 * 2^(-35+1) + ( 1^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = 1 
assign u[4'b1001] [35] = 21'h 0007FF;  // +1.9999999999854481 = 2^36 * ln( 1 +  1 * 2^(-36+1) + ( 1^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = 1 
assign u[4'b1001] [36] = 21'h 0007FF;  // +1.9999999999927240 = 2^37 * ln( 1 +  1 * 2^(-37+1) + ( 1^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = 1 
assign u[4'b1001] [37] = 21'h 0007FF;  // +1.9999999999963620 = 2^38 * ln( 1 +  1 * 2^(-38+1) + ( 1^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = 1 
assign u[4'b1001] [38] = 21'h 0007FF;  // +1.9999999999981810 = 2^39 * ln( 1 +  1 * 2^(-39+1) + ( 1^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = 1 
assign u[4'b1001] [39] = 21'h 0007FF;  // +1.9999999999990905 = 2^40 * ln( 1 +  1 * 2^(-40+1) + ( 1^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = 1 
assign u[4'b1001] [40] = 21'h 0007FF;  // +1.9999999999995453 = 2^41 * ln( 1 +  1 * 2^(-41+1) + ( 1^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = 1 
assign u[4'b1001] [41] = 21'h 0007FF;  // +1.9999999999997726 = 2^42 * ln( 1 +  1 * 2^(-42+1) + ( 1^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = 1 
assign u[4'b1001] [42] = 21'h 0007FF;  // +1.9999999999998863 = 2^43 * ln( 1 +  1 * 2^(-43+1) + ( 1^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = 1 
assign u[4'b1001] [43] = 21'h 0007FF;  // +1.9999999999999432 = 2^44 * ln( 1 +  1 * 2^(-44+1) + ( 1^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = 1 
assign u[4'b1001] [44] = 21'h 0007FF;  // +1.9999999999999716 = 2^45 * ln( 1 +  1 * 2^(-45+1) + ( 1^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = 1 
assign u[4'b1001] [45] = 21'h 0007FF;  // +1.9999999999999858 = 2^46 * ln( 1 +  1 * 2^(-46+1) + ( 1^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = 1 
assign u[4'b1001] [46] = 21'h 0007FF;  // +1.9999999999999929 = 2^47 * ln( 1 +  1 * 2^(-47+1) + ( 1^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = 1 
assign u[4'b1001] [47] = 21'h 0007FF;  // +1.9999999999999964 = 2^48 * ln( 1 +  1 * 2^(-48+1) + ( 1^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = 1 
assign u[4'b1001] [48] = 21'h 0007FF;  // +1.9999999999999982 = 2^49 * ln( 1 +  1 * 2^(-49+1) + ( 1^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = 1 
assign u[4'b1001] [49] = 21'h 0007FF;  // +1.9999999999999991 = 2^50 * ln( 1 +  1 * 2^(-50+1) + ( 1^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = 1 
assign u[4'b1001] [50] = 21'h 0007FF;  // +1.9999999999999996 = 2^51 * ln( 1 +  1 * 2^(-51+1) + ( 1^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = 1 
assign u[4'b1001] [51] = 21'h 0007FF;  // +1.9999999999999998 = 2^52 * ln( 1 +  1 * 2^(-52+1) + ( 1^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = 1 
assign u[4'b1001] [52] = 21'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  1 * 2^(-53+1) + ( 1^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = 1 
assign u[4'b1001] [53] = 21'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  1 * 2^(-54+1) + ( 1^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = 1 
assign u[4'b1001] [54] = 21'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  1 * 2^(-55+1) + ( 1^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = 1 
assign u[4'b1001] [55] = 21'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  1 * 2^(-56+1) + ( 1^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = 1 
assign u[4'b1001] [56] = 21'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  1 * 2^(-57+1) + ( 1^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = 1 
assign u[4'b1001] [57] = 21'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  1 * 2^(-58+1) + ( 1^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = 1 
assign u[4'b1001] [58] = 21'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  1 * 2^(-59+1) + ( 1^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = 1 
assign u[4'b1001] [59] = 21'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  1 * 2^(-60+1) + ( 1^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = 1 
assign u[4'b1001] [60] = 21'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  1 * 2^(-61+1) + ( 1^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = 1 
assign u[4'b1001] [61] = 21'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  1 * 2^(-62+1) + ( 1^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = 1 
assign u[4'b1001] [62] = 21'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  1 * 2^(-63+1) + ( 1^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = 1 
assign u[4'b1001] [63] = 21'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  1 * 2^(-64+1) + ( 1^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = 1 
assign u[4'b1010] [00] = 21'h 000000;  // +0.0000000000000000 = 2^ 1 * ln( 1 +  0 * 2^(- 1+1) + ( 0^2+ 0^2) * 2^(-2* 1) )   n =  1   d_n = -0 
assign u[4'b1010] [01] = 21'h 000000;  // +0.0000000000000000 = 2^ 2 * ln( 1 +  0 * 2^(- 2+1) + ( 0^2+ 0^2) * 2^(-2* 2) )   n =  2   d_n = -0 
assign u[4'b1010] [02] = 21'h 000000;  // +0.0000000000000000 = 2^ 3 * ln( 1 +  0 * 2^(- 3+1) + ( 0^2+ 0^2) * 2^(-2* 3) )   n =  3   d_n = -0 
assign u[4'b1010] [03] = 21'h 000000;  // +0.0000000000000000 = 2^ 4 * ln( 1 +  0 * 2^(- 4+1) + ( 0^2+ 0^2) * 2^(-2* 4) )   n =  4   d_n = -0 
assign u[4'b1010] [04] = 21'h 000000;  // +0.0000000000000000 = 2^ 5 * ln( 1 +  0 * 2^(- 5+1) + ( 0^2+ 0^2) * 2^(-2* 5) )   n =  5   d_n = -0 
assign u[4'b1010] [05] = 21'h 000000;  // +0.0000000000000000 = 2^ 6 * ln( 1 +  0 * 2^(- 6+1) + ( 0^2+ 0^2) * 2^(-2* 6) )   n =  6   d_n = -0 
assign u[4'b1010] [06] = 21'h 000000;  // +0.0000000000000000 = 2^ 7 * ln( 1 +  0 * 2^(- 7+1) + ( 0^2+ 0^2) * 2^(-2* 7) )   n =  7   d_n = -0 
assign u[4'b1010] [07] = 21'h 000000;  // +0.0000000000000000 = 2^ 8 * ln( 1 +  0 * 2^(- 8+1) + ( 0^2+ 0^2) * 2^(-2* 8) )   n =  8   d_n = -0 
assign u[4'b1010] [08] = 21'h 000000;  // +0.0000000000000000 = 2^ 9 * ln( 1 +  0 * 2^(- 9+1) + ( 0^2+ 0^2) * 2^(-2* 9) )   n =  9   d_n = -0 
assign u[4'b1010] [09] = 21'h 000000;  // +0.0000000000000000 = 2^10 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = -0 
assign u[4'b1010] [10] = 21'h 000000;  // +0.0000000000000000 = 2^11 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = -0 
assign u[4'b1010] [11] = 21'h 000000;  // +0.0000000000000000 = 2^12 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = -0 
assign u[4'b1010] [12] = 21'h 000000;  // +0.0000000000000000 = 2^13 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = -0 
assign u[4'b1010] [13] = 21'h 000000;  // +0.0000000000000000 = 2^14 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = -0 
assign u[4'b1010] [14] = 21'h 000000;  // +0.0000000000000000 = 2^15 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = -0 
assign u[4'b1010] [15] = 21'h 000000;  // +0.0000000000000000 = 2^16 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = -0 
assign u[4'b1010] [16] = 21'h 000000;  // +0.0000000000000000 = 2^17 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = -0 
assign u[4'b1010] [17] = 21'h 000000;  // +0.0000000000000000 = 2^18 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = -0 
assign u[4'b1010] [18] = 21'h 000000;  // +0.0000000000000000 = 2^19 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = -0 
assign u[4'b1010] [19] = 21'h 000000;  // +0.0000000000000000 = 2^20 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = -0 
assign u[4'b1010] [20] = 21'h 000000;  // +0.0000000000000000 = 2^21 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = -0 
assign u[4'b1010] [21] = 21'h 000000;  // +0.0000000000000000 = 2^22 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = -0 
assign u[4'b1010] [22] = 21'h 000000;  // +0.0000000000000000 = 2^23 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = -0 
assign u[4'b1010] [23] = 21'h 000000;  // +0.0000000000000000 = 2^24 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = -0 
assign u[4'b1010] [24] = 21'h 000000;  // +0.0000000000000000 = 2^25 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = -0 
assign u[4'b1010] [25] = 21'h 000000;  // +0.0000000000000000 = 2^26 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = -0 
assign u[4'b1010] [26] = 21'h 000000;  // +0.0000000000000000 = 2^27 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = -0 
assign u[4'b1010] [27] = 21'h 000000;  // +0.0000000000000000 = 2^28 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = -0 
assign u[4'b1010] [28] = 21'h 000000;  // +0.0000000000000000 = 2^29 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = -0 
assign u[4'b1010] [29] = 21'h 000000;  // +0.0000000000000000 = 2^30 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = -0 
assign u[4'b1010] [30] = 21'h 000000;  // +0.0000000000000000 = 2^31 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = -0 
assign u[4'b1010] [31] = 21'h 000000;  // +0.0000000000000000 = 2^32 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = -0 
assign u[4'b1010] [32] = 21'h 000000;  // +0.0000000000000000 = 2^33 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = -0 
assign u[4'b1010] [33] = 21'h 000000;  // +0.0000000000000000 = 2^34 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = -0 
assign u[4'b1010] [34] = 21'h 000000;  // +0.0000000000000000 = 2^35 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = -0 
assign u[4'b1010] [35] = 21'h 000000;  // +0.0000000000000000 = 2^36 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = -0 
assign u[4'b1010] [36] = 21'h 000000;  // +0.0000000000000000 = 2^37 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = -0 
assign u[4'b1010] [37] = 21'h 000000;  // +0.0000000000000000 = 2^38 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = -0 
assign u[4'b1010] [38] = 21'h 000000;  // +0.0000000000000000 = 2^39 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = -0 
assign u[4'b1010] [39] = 21'h 000000;  // +0.0000000000000000 = 2^40 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = -0 
assign u[4'b1010] [40] = 21'h 000000;  // +0.0000000000000000 = 2^41 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = -0 
assign u[4'b1010] [41] = 21'h 000000;  // +0.0000000000000000 = 2^42 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = -0 
assign u[4'b1010] [42] = 21'h 000000;  // +0.0000000000000000 = 2^43 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = -0 
assign u[4'b1010] [43] = 21'h 000000;  // +0.0000000000000000 = 2^44 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = -0 
assign u[4'b1010] [44] = 21'h 000000;  // +0.0000000000000000 = 2^45 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = -0 
assign u[4'b1010] [45] = 21'h 000000;  // +0.0000000000000000 = 2^46 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = -0 
assign u[4'b1010] [46] = 21'h 000000;  // +0.0000000000000000 = 2^47 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = -0 
assign u[4'b1010] [47] = 21'h 000000;  // +0.0000000000000000 = 2^48 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = -0 
assign u[4'b1010] [48] = 21'h 000000;  // +0.0000000000000000 = 2^49 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = -0 
assign u[4'b1010] [49] = 21'h 000000;  // +0.0000000000000000 = 2^50 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = -0 
assign u[4'b1010] [50] = 21'h 000000;  // +0.0000000000000000 = 2^51 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = -0 
assign u[4'b1010] [51] = 21'h 000000;  // +0.0000000000000000 = 2^52 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = -0 
assign u[4'b1010] [52] = 21'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = -0 
assign u[4'b1010] [53] = 21'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = -0 
assign u[4'b1010] [54] = 21'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = -0 
assign u[4'b1010] [55] = 21'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = -0 
assign u[4'b1010] [56] = 21'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = -0 
assign u[4'b1010] [57] = 21'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = -0 
assign u[4'b1010] [58] = 21'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = -0 
assign u[4'b1010] [59] = 21'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = -0 
assign u[4'b1010] [60] = 21'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = -0 
assign u[4'b1010] [61] = 21'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = -0 
assign u[4'b1010] [62] = 21'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = -0 
assign u[4'b1010] [63] = 21'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = -0 
assign u[4'b1011] [00] = 21'h 1FF4E8;  // -2.7725887222397811 = 2^ 1 * ln( 1 + -1 * 2^(- 1+1) + (-1^2+ 0^2) * 2^(-2* 1) )   n =  1   d_n = -1 
assign u[4'b1011] [01] = 21'h 1FF6CB;  // -2.3014565796142472 = 2^ 2 * ln( 1 + -1 * 2^(- 2+1) + (-1^2+ 0^2) * 2^(-2* 2) )   n =  2   d_n = -1 
assign u[4'b1011] [02] = 21'h 1FF774;  // -2.1365022819923620 = 2^ 3 * ln( 1 + -1 * 2^(- 3+1) + (-1^2+ 0^2) * 2^(-2* 3) )   n =  3   d_n = -1 
assign u[4'b1011] [03] = 21'h 1FF7BD;  // -2.0652326764022777 = 2^ 4 * ln( 1 + -1 * 2^(- 4+1) + (-1^2+ 0^2) * 2^(-2* 4) )   n =  4   d_n = -1 
assign u[4'b1011] [04] = 21'h 1FF7DF;  // -2.0319166921331391 = 2^ 5 * ln( 1 + -1 * 2^(- 5+1) + (-1^2+ 0^2) * 2^(-2* 5) )   n =  5   d_n = -1 
assign u[4'b1011] [05] = 21'h 1FF7EF;  // -2.0157896919218135 = 2^ 6 * ln( 1 + -1 * 2^(- 6+1) + (-1^2+ 0^2) * 2^(-2* 6) )   n =  6   d_n = -1 
assign u[4'b1011] [06] = 21'h 1FF7F7;  // -2.0078534300226285 = 2^ 7 * ln( 1 + -1 * 2^(- 7+1) + (-1^2+ 0^2) * 2^(-2* 7) )   n =  7   d_n = -1 
assign u[4'b1011] [07] = 21'h 1FF7FB;  // -2.0039164524218003 = 2^ 8 * ln( 1 + -1 * 2^(- 8+1) + (-1^2+ 0^2) * 2^(-2* 8) )   n =  8   d_n = -1 
assign u[4'b1011] [08] = 21'h 1FF7FD;  // -2.0019556718626310 = 2^ 9 * ln( 1 + -1 * 2^(- 9+1) + (-1^2+ 0^2) * 2^(-2* 9) )   n =  9   d_n = -1 
assign u[4'b1011] [09] = 21'h 1FF7FE;  // -2.0009771987489029 = 2^10 * ln( 1 + -1 * 2^(-10+1) + (-1^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = -1 
assign u[4'b1011] [10] = 21'h 1FF7FF;  // -2.0004884402539500 = 2^11 * ln( 1 + -1 * 2^(-11+1) + (-1^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = -1 
assign u[4'b1011] [11] = 21'h 1FF7FF;  // -2.0002441803687074 = 2^12 * ln( 1 + -1 * 2^(-12+1) + (-1^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = -1 
assign u[4'b1011] [12] = 21'h 1FF7FF;  // -2.0001220802475173 = 2^13 * ln( 1 + -1 * 2^(-13+1) + (-1^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = -1 
assign u[4'b1011] [13] = 21'h 1FF7FF;  // -2.0000610376398904 = 2^14 * ln( 1 + -1 * 2^(-14+1) + (-1^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = -1 
assign u[4'b1011] [14] = 21'h 1FF7FF;  // -2.0000305181990208 = 2^15 * ln( 1 + -1 * 2^(-15+1) + (-1^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = -1 
assign u[4'b1011] [15] = 21'h 1FF7FF;  // -2.0000152589442846 = 2^16 * ln( 1 + -1 * 2^(-16+1) + (-1^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = -1 
assign u[4'b1011] [16] = 21'h 1FF7FF;  // -2.0000076294333367 = 2^17 * ln( 1 + -1 * 2^(-17+1) + (-1^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = -1 
assign u[4'b1011] [17] = 21'h 1FF7FF;  // -2.0000038147069668 = 2^18 * ln( 1 + -1 * 2^(-18+1) + (-1^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = -1 
assign u[4'b1011] [18] = 21'h 1FF7FF;  // -2.0000019073510580 = 2^19 * ln( 1 + -1 * 2^(-19+1) + (-1^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = -1 
assign u[4'b1011] [19] = 21'h 1FF7FF;  // -2.0000009536749226 = 2^20 * ln( 1 + -1 * 2^(-20+1) + (-1^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = -1 
assign u[4'b1011] [20] = 21'h 1FF7FF;  // -2.0000004768373096 = 2^21 * ln( 1 + -1 * 2^(-21+1) + (-1^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = -1 
assign u[4'b1011] [21] = 21'h 1FF7FF;  // -2.0000002384186168 = 2^22 * ln( 1 + -1 * 2^(-22+1) + (-1^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = -1 
assign u[4'b1011] [22] = 21'h 1FF7FF;  // -2.0000001192092989 = 2^23 * ln( 1 + -1 * 2^(-23+1) + (-1^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = -1 
assign u[4'b1011] [23] = 21'h 1FF7FF;  // -2.0000000596046470 = 2^24 * ln( 1 + -1 * 2^(-24+1) + (-1^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = -1 
assign u[4'b1011] [24] = 21'h 1FF7FF;  // -2.0000000298023228 = 2^25 * ln( 1 + -1 * 2^(-25+1) + (-1^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = -1 
assign u[4'b1011] [25] = 21'h 1FF7FF;  // -2.0000000149011612 = 2^26 * ln( 1 + -1 * 2^(-26+1) + (-1^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = -1 
assign u[4'b1011] [26] = 21'h 1FF7FF;  // -2.0000000074505806 = 2^27 * ln( 1 + -1 * 2^(-27+1) + (-1^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = -1 
assign u[4'b1011] [27] = 21'h 1FF7FF;  // -2.0000000037252903 = 2^28 * ln( 1 + -1 * 2^(-28+1) + (-1^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = -1 
assign u[4'b1011] [28] = 21'h 1FF7FF;  // -2.0000000018626451 = 2^29 * ln( 1 + -1 * 2^(-29+1) + (-1^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = -1 
assign u[4'b1011] [29] = 21'h 1FF7FF;  // -2.0000000009313226 = 2^30 * ln( 1 + -1 * 2^(-30+1) + (-1^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = -1 
assign u[4'b1011] [30] = 21'h 1FF7FF;  // -2.0000000004656613 = 2^31 * ln( 1 + -1 * 2^(-31+1) + (-1^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = -1 
assign u[4'b1011] [31] = 21'h 1FF7FF;  // -2.0000000002328306 = 2^32 * ln( 1 + -1 * 2^(-32+1) + (-1^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = -1 
assign u[4'b1011] [32] = 21'h 1FF7FF;  // -2.0000000001164153 = 2^33 * ln( 1 + -1 * 2^(-33+1) + (-1^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = -1 
assign u[4'b1011] [33] = 21'h 1FF7FF;  // -2.0000000000582077 = 2^34 * ln( 1 + -1 * 2^(-34+1) + (-1^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = -1 
assign u[4'b1011] [34] = 21'h 1FF7FF;  // -2.0000000000291038 = 2^35 * ln( 1 + -1 * 2^(-35+1) + (-1^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = -1 
assign u[4'b1011] [35] = 21'h 1FF7FF;  // -2.0000000000145519 = 2^36 * ln( 1 + -1 * 2^(-36+1) + (-1^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = -1 
assign u[4'b1011] [36] = 21'h 1FF7FF;  // -2.0000000000072760 = 2^37 * ln( 1 + -1 * 2^(-37+1) + (-1^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = -1 
assign u[4'b1011] [37] = 21'h 1FF7FF;  // -2.0000000000036380 = 2^38 * ln( 1 + -1 * 2^(-38+1) + (-1^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = -1 
assign u[4'b1011] [38] = 21'h 1FF7FF;  // -2.0000000000018190 = 2^39 * ln( 1 + -1 * 2^(-39+1) + (-1^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = -1 
assign u[4'b1011] [39] = 21'h 1FF7FF;  // -2.0000000000009095 = 2^40 * ln( 1 + -1 * 2^(-40+1) + (-1^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = -1 
assign u[4'b1011] [40] = 21'h 1FF7FF;  // -2.0000000000004547 = 2^41 * ln( 1 + -1 * 2^(-41+1) + (-1^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = -1 
assign u[4'b1011] [41] = 21'h 1FF7FF;  // -2.0000000000002274 = 2^42 * ln( 1 + -1 * 2^(-42+1) + (-1^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = -1 
assign u[4'b1011] [42] = 21'h 1FF800;  // -2.0000000000001137 = 2^43 * ln( 1 + -1 * 2^(-43+1) + (-1^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = -1 
assign u[4'b1011] [43] = 21'h 1FF800;  // -2.0000000000000568 = 2^44 * ln( 1 + -1 * 2^(-44+1) + (-1^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = -1 
assign u[4'b1011] [44] = 21'h 1FF800;  // -2.0000000000000284 = 2^45 * ln( 1 + -1 * 2^(-45+1) + (-1^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = -1 
assign u[4'b1011] [45] = 21'h 1FF800;  // -2.0000000000000142 = 2^46 * ln( 1 + -1 * 2^(-46+1) + (-1^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = -1 
assign u[4'b1011] [46] = 21'h 1FF800;  // -2.0000000000000071 = 2^47 * ln( 1 + -1 * 2^(-47+1) + (-1^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = -1 
assign u[4'b1011] [47] = 21'h 1FF800;  // -2.0000000000000036 = 2^48 * ln( 1 + -1 * 2^(-48+1) + (-1^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = -1 
assign u[4'b1011] [48] = 21'h 1FF800;  // -2.0000000000000018 = 2^49 * ln( 1 + -1 * 2^(-49+1) + (-1^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = -1 
assign u[4'b1011] [49] = 21'h 1FF800;  // -2.0000000000000009 = 2^50 * ln( 1 + -1 * 2^(-50+1) + (-1^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = -1 
assign u[4'b1011] [50] = 21'h 1FF800;  // -2.0000000000000004 = 2^51 * ln( 1 + -1 * 2^(-51+1) + (-1^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = -1 
assign u[4'b1011] [51] = 21'h 1FF800;  // -2.0000000000000004 = 2^52 * ln( 1 + -1 * 2^(-52+1) + (-1^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = -1 
assign u[4'b1011] [52] = 21'h 1FF800;  // -2.0000000000000000 = 2^53 * ln( 1 + -1 * 2^(-53+1) + (-1^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = -1 
assign u[4'b1011] [53] = 21'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 + -1 * 2^(-54+1) + (-1^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = -1 
assign u[4'b1011] [54] = 21'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 + -1 * 2^(-55+1) + (-1^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = -1 
assign u[4'b1011] [55] = 21'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 + -1 * 2^(-56+1) + (-1^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = -1 
assign u[4'b1011] [56] = 21'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 + -1 * 2^(-57+1) + (-1^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = -1 
assign u[4'b1011] [57] = 21'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 + -1 * 2^(-58+1) + (-1^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = -1 
assign u[4'b1011] [58] = 21'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 + -1 * 2^(-59+1) + (-1^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = -1 
assign u[4'b1011] [59] = 21'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 + -1 * 2^(-60+1) + (-1^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = -1 
assign u[4'b1011] [60] = 21'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 + -1 * 2^(-61+1) + (-1^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = -1 
assign u[4'b1011] [61] = 21'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 + -1 * 2^(-62+1) + (-1^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = -1 
assign u[4'b1011] [62] = 21'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 + -1 * 2^(-63+1) + (-1^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = -1 
assign u[4'b1011] [63] = 21'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 + -1 * 2^(-64+1) + (-1^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = -1 
assign u[4'b1100] [00] = 21'h 0001C8;  // +0.4462871026284197 = 2^ 1 * ln( 1 +  0 * 2^(- 1+1) + ( 0^2+-1^2) * 2^(-2* 1) )   n =  1   d_n = -0-1i 
assign u[4'b1100] [01] = 21'h 0000F8;  // +0.2424984872657394 = 2^ 2 * ln( 1 +  0 * 2^(- 2+1) + ( 0^2+-1^2) * 2^(-2* 2) )   n =  2   d_n = -0-1i 
assign u[4'b1100] [02] = 21'h 00007F;  // +0.1240334922877210 = 2^ 3 * ln( 1 +  0 * 2^(- 3+1) + ( 0^2+-1^2) * 2^(-2* 3) )   n =  3   d_n = -0-1i 
assign u[4'b1100] [03] = 21'h 00003F;  // +0.0623782466505195 = 2^ 4 * ln( 1 +  0 * 2^(- 4+1) + ( 0^2+-1^2) * 2^(-2* 4) )   n =  4   d_n = -0-1i 
assign u[4'b1100] [04] = 21'h 00001F;  // +0.0312347511377731 = 2^ 5 * ln( 1 +  0 * 2^(- 5+1) + ( 0^2+-1^2) * 2^(-2* 5) )   n =  5   d_n = -0-1i 
assign u[4'b1100] [05] = 21'h 00000F;  // +0.0156230929617406 = 2^ 6 * ln( 1 +  0 * 2^(- 6+1) + ( 0^2+-1^2) * 2^(-2* 6) )   n =  6   d_n = -0-1i 
assign u[4'b1100] [06] = 21'h 000007;  // +0.0078122615911219 = 2^ 7 * ln( 1 +  0 * 2^(- 7+1) + ( 0^2+-1^2) * 2^(-2* 7) )   n =  7   d_n = -0-1i 
assign u[4'b1100] [07] = 21'h 000003;  // +0.0039062201979808 = 2^ 8 * ln( 1 +  0 * 2^(- 8+1) + ( 0^2+-1^2) * 2^(-2* 8) )   n =  8   d_n = -0-1i 
assign u[4'b1100] [08] = 21'h 000001;  // +0.0019531212747156 = 2^ 9 * ln( 1 +  0 * 2^(- 9+1) + ( 0^2+-1^2) * 2^(-2* 9) )   n =  9   d_n = -0-1i 
assign u[4'b1100] [09] = 21'h 000000;  // +0.0009765620343389 = 2^10 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+-1^2) * 2^(-2*10) )   n = 10   d_n = -0-1i 
assign u[4'b1100] [10] = 21'h 000000;  // +0.0004882811917923 = 2^11 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+-1^2) * 2^(-2*11) )   n = 11   d_n = -0-1i 
assign u[4'b1100] [11] = 21'h 000000;  // +0.0002441406177240 = 2^12 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+-1^2) * 2^(-2*12) )   n = 12   d_n = -0-1i 
assign u[4'b1100] [12] = 21'h 000000;  // +0.0001220703120453 = 2^13 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+-1^2) * 2^(-2*13) )   n = 13   d_n = -0-1i 
assign u[4'b1100] [13] = 21'h 000000;  // +0.0000610351561932 = 2^14 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+-1^2) * 2^(-2*14) )   n = 14   d_n = -0-1i 
assign u[4'b1100] [14] = 21'h 000000;  // +0.0000305175781179 = 2^15 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+-1^2) * 2^(-2*15) )   n = 15   d_n = -0-1i 
assign u[4'b1100] [15] = 21'h 000000;  // +0.0000152587890616 = 2^16 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+-1^2) * 2^(-2*16) )   n = 16   d_n = -0-1i 
assign u[4'b1100] [16] = 21'h 000000;  // +0.0000076293945311 = 2^17 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+-1^2) * 2^(-2*17) )   n = 17   d_n = -0-1i 
assign u[4'b1100] [17] = 21'h 000000;  // +0.0000038146972656 = 2^18 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+-1^2) * 2^(-2*18) )   n = 18   d_n = -0-1i 
assign u[4'b1100] [18] = 21'h 000000;  // +0.0000019073486328 = 2^19 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+-1^2) * 2^(-2*19) )   n = 19   d_n = -0-1i 
assign u[4'b1100] [19] = 21'h 000000;  // +0.0000009536743164 = 2^20 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+-1^2) * 2^(-2*20) )   n = 20   d_n = -0-1i 
assign u[4'b1100] [20] = 21'h 000000;  // +0.0000004768371582 = 2^21 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+-1^2) * 2^(-2*21) )   n = 21   d_n = -0-1i 
assign u[4'b1100] [21] = 21'h 000000;  // +0.0000002384185791 = 2^22 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+-1^2) * 2^(-2*22) )   n = 22   d_n = -0-1i 
assign u[4'b1100] [22] = 21'h 000000;  // +0.0000001192092896 = 2^23 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+-1^2) * 2^(-2*23) )   n = 23   d_n = -0-1i 
assign u[4'b1100] [23] = 21'h 000000;  // +0.0000000596046448 = 2^24 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+-1^2) * 2^(-2*24) )   n = 24   d_n = -0-1i 
assign u[4'b1100] [24] = 21'h 000000;  // +0.0000000298023224 = 2^25 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+-1^2) * 2^(-2*25) )   n = 25   d_n = -0-1i 
assign u[4'b1100] [25] = 21'h 000000;  // +0.0000000000000000 = 2^26 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+-1^2) * 2^(-2*26) )   n = 26   d_n = -0-1i 
assign u[4'b1100] [26] = 21'h 000000;  // +0.0000000000000000 = 2^27 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+-1^2) * 2^(-2*27) )   n = 27   d_n = -0-1i 
assign u[4'b1100] [27] = 21'h 000000;  // +0.0000000000000000 = 2^28 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+-1^2) * 2^(-2*28) )   n = 28   d_n = -0-1i 
assign u[4'b1100] [28] = 21'h 000000;  // +0.0000000000000000 = 2^29 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+-1^2) * 2^(-2*29) )   n = 29   d_n = -0-1i 
assign u[4'b1100] [29] = 21'h 000000;  // +0.0000000000000000 = 2^30 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+-1^2) * 2^(-2*30) )   n = 30   d_n = -0-1i 
assign u[4'b1100] [30] = 21'h 000000;  // +0.0000000000000000 = 2^31 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+-1^2) * 2^(-2*31) )   n = 31   d_n = -0-1i 
assign u[4'b1100] [31] = 21'h 000000;  // +0.0000000000000000 = 2^32 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+-1^2) * 2^(-2*32) )   n = 32   d_n = -0-1i 
assign u[4'b1100] [32] = 21'h 000000;  // +0.0000000000000000 = 2^33 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+-1^2) * 2^(-2*33) )   n = 33   d_n = -0-1i 
assign u[4'b1100] [33] = 21'h 000000;  // +0.0000000000000000 = 2^34 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+-1^2) * 2^(-2*34) )   n = 34   d_n = -0-1i 
assign u[4'b1100] [34] = 21'h 000000;  // +0.0000000000000000 = 2^35 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+-1^2) * 2^(-2*35) )   n = 35   d_n = -0-1i 
assign u[4'b1100] [35] = 21'h 000000;  // +0.0000000000000000 = 2^36 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+-1^2) * 2^(-2*36) )   n = 36   d_n = -0-1i 
assign u[4'b1100] [36] = 21'h 000000;  // +0.0000000000000000 = 2^37 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+-1^2) * 2^(-2*37) )   n = 37   d_n = -0-1i 
assign u[4'b1100] [37] = 21'h 000000;  // +0.0000000000000000 = 2^38 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+-1^2) * 2^(-2*38) )   n = 38   d_n = -0-1i 
assign u[4'b1100] [38] = 21'h 000000;  // +0.0000000000000000 = 2^39 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+-1^2) * 2^(-2*39) )   n = 39   d_n = -0-1i 
assign u[4'b1100] [39] = 21'h 000000;  // +0.0000000000000000 = 2^40 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+-1^2) * 2^(-2*40) )   n = 40   d_n = -0-1i 
assign u[4'b1100] [40] = 21'h 000000;  // +0.0000000000000000 = 2^41 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+-1^2) * 2^(-2*41) )   n = 41   d_n = -0-1i 
assign u[4'b1100] [41] = 21'h 000000;  // +0.0000000000000000 = 2^42 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+-1^2) * 2^(-2*42) )   n = 42   d_n = -0-1i 
assign u[4'b1100] [42] = 21'h 000000;  // +0.0000000000000000 = 2^43 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+-1^2) * 2^(-2*43) )   n = 43   d_n = -0-1i 
assign u[4'b1100] [43] = 21'h 000000;  // +0.0000000000000000 = 2^44 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+-1^2) * 2^(-2*44) )   n = 44   d_n = -0-1i 
assign u[4'b1100] [44] = 21'h 000000;  // +0.0000000000000000 = 2^45 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+-1^2) * 2^(-2*45) )   n = 45   d_n = -0-1i 
assign u[4'b1100] [45] = 21'h 000000;  // +0.0000000000000000 = 2^46 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+-1^2) * 2^(-2*46) )   n = 46   d_n = -0-1i 
assign u[4'b1100] [46] = 21'h 000000;  // +0.0000000000000000 = 2^47 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+-1^2) * 2^(-2*47) )   n = 47   d_n = -0-1i 
assign u[4'b1100] [47] = 21'h 000000;  // +0.0000000000000000 = 2^48 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+-1^2) * 2^(-2*48) )   n = 48   d_n = -0-1i 
assign u[4'b1100] [48] = 21'h 000000;  // +0.0000000000000000 = 2^49 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+-1^2) * 2^(-2*49) )   n = 49   d_n = -0-1i 
assign u[4'b1100] [49] = 21'h 000000;  // +0.0000000000000000 = 2^50 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+-1^2) * 2^(-2*50) )   n = 50   d_n = -0-1i 
assign u[4'b1100] [50] = 21'h 000000;  // +0.0000000000000000 = 2^51 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+-1^2) * 2^(-2*51) )   n = 51   d_n = -0-1i 
assign u[4'b1100] [51] = 21'h 000000;  // +0.0000000000000000 = 2^52 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+-1^2) * 2^(-2*52) )   n = 52   d_n = -0-1i 
assign u[4'b1100] [52] = 21'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+-1^2) * 2^(-2*53) )   n = 53   d_n = -0-1i 
assign u[4'b1100] [53] = 21'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+-1^2) * 2^(-2*54) )   n = 54   d_n = -0-1i 
assign u[4'b1100] [54] = 21'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+-1^2) * 2^(-2*55) )   n = 55   d_n = -0-1i 
assign u[4'b1100] [55] = 21'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+-1^2) * 2^(-2*56) )   n = 56   d_n = -0-1i 
assign u[4'b1100] [56] = 21'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+-1^2) * 2^(-2*57) )   n = 57   d_n = -0-1i 
assign u[4'b1100] [57] = 21'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+-1^2) * 2^(-2*58) )   n = 58   d_n = -0-1i 
assign u[4'b1100] [58] = 21'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+-1^2) * 2^(-2*59) )   n = 59   d_n = -0-1i 
assign u[4'b1100] [59] = 21'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+-1^2) * 2^(-2*60) )   n = 60   d_n = -0-1i 
assign u[4'b1100] [60] = 21'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+-1^2) * 2^(-2*61) )   n = 61   d_n = -0-1i 
assign u[4'b1100] [61] = 21'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+-1^2) * 2^(-2*62) )   n = 62   d_n = -0-1i 
assign u[4'b1100] [62] = 21'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+-1^2) * 2^(-2*63) )   n = 63   d_n = -0-1i 
assign u[4'b1100] [63] = 21'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+-1^2) * 2^(-2*64) )   n = 64   d_n = -0-1i 
assign u[4'b1101] [00] = 21'h 000754;  // +1.8325814637483104 = 2^ 1 * ln( 1 +  1 * 2^(- 1+1) + ( 1^2+-1^2) * 2^(-2* 1) )   n =  1   d_n = 1-1i 
assign u[4'b1101] [01] = 21'h 0007C4;  // +1.9420312631268026 = 2^ 2 * ln( 1 +  1 * 2^(- 2+1) + ( 1^2+-1^2) * 2^(-2* 2) )   n =  2   d_n = 1-1i 
assign u[4'b1101] [02] = 21'h 0007EE;  // +1.9826893112366513 = 2^ 3 * ln( 1 +  1 * 2^(- 3+1) + ( 1^2+-1^2) * 2^(-2* 3) )   n =  3   d_n = 1-1i 
assign u[4'b1101] [03] = 21'h 0007FB;  // +1.9952556560153185 = 2^ 4 * ln( 1 +  1 * 2^(- 4+1) + ( 1^2+-1^2) * 2^(-2* 4) )   n =  4   d_n = 1-1i 
assign u[4'b1101] [04] = 21'h 0007FE;  // +1.9987574279595595 = 2^ 5 * ln( 1 +  1 * 2^(- 5+1) + ( 1^2+-1^2) * 2^(-2* 5) )   n =  5   d_n = 1-1i 
assign u[4'b1101] [05] = 21'h 0007FF;  // +1.9996820132261188 = 2^ 6 * ln( 1 +  1 * 2^(- 6+1) + ( 1^2+-1^2) * 2^(-2* 6) )   n =  6   d_n = 1-1i 
assign u[4'b1101] [06] = 21'h 0007FF;  // +1.9999195675060046 = 2^ 7 * ln( 1 +  1 * 2^(- 7+1) + ( 1^2+-1^2) * 2^(-2* 7) )   n =  7   d_n = 1-1i 
assign u[4'b1101] [07] = 21'h 0007FF;  // +1.9999797737846823 = 2^ 8 * ln( 1 +  1 * 2^(- 8+1) + ( 1^2+-1^2) * 2^(-2* 8) )   n =  8   d_n = 1-1i 
assign u[4'b1101] [08] = 21'h 0007FF;  // +1.9999949286148679 = 2^ 9 * ln( 1 +  1 * 2^(- 9+1) + ( 1^2+-1^2) * 2^(-2* 9) )   n =  9   d_n = 1-1i 
assign u[4'b1101] [09] = 21'h 0007FF;  // +1.9999987302952080 = 2^10 * ln( 1 +  1 * 2^(-10+1) + ( 1^2+-1^2) * 2^(-2*10) )   n = 10   d_n = 1-1i 
assign u[4'b1101] [10] = 21'h 0007FF;  // +1.9999996823413151 = 2^11 * ln( 1 +  1 * 2^(-11+1) + ( 1^2+-1^2) * 2^(-2*11) )   n = 11   d_n = 1-1i 
assign u[4'b1101] [11] = 21'h 0007FF;  // +1.9999999205562393 = 2^12 * ln( 1 +  1 * 2^(-12+1) + ( 1^2+-1^2) * 2^(-2*12) )   n = 12   d_n = 1-1i 
assign u[4'b1101] [12] = 21'h 0007FF;  // +1.9999999801340587 = 2^13 * ln( 1 +  1 * 2^(-13+1) + ( 1^2+-1^2) * 2^(-2*13) )   n = 13   d_n = 1-1i 
assign u[4'b1101] [13] = 21'h 0007FF;  // +1.9999999950332306 = 2^14 * ln( 1 +  1 * 2^(-14+1) + ( 1^2+-1^2) * 2^(-2*14) )   n = 14   d_n = 1-1i 
assign u[4'b1101] [14] = 21'h 0007FF;  // +1.9999999987582722 = 2^15 * ln( 1 +  1 * 2^(-15+1) + ( 1^2+-1^2) * 2^(-2*15) )   n = 15   d_n = 1-1i 
assign u[4'b1101] [15] = 21'h 0007FF;  // +1.9999999996895637 = 2^16 * ln( 1 +  1 * 2^(-16+1) + ( 1^2+-1^2) * 2^(-2*16) )   n = 16   d_n = 1-1i 
assign u[4'b1101] [16] = 21'h 0007FF;  // +1.9999999999223903 = 2^17 * ln( 1 +  1 * 2^(-17+1) + ( 1^2+-1^2) * 2^(-2*17) )   n = 17   d_n = 1-1i 
assign u[4'b1101] [17] = 21'h 0007FF;  // +1.9999999999951494 = 2^18 * ln( 1 +  1 * 2^(-18+1) + ( 1^2+-1^2) * 2^(-2*18) )   n = 18   d_n = 1-1i 
assign u[4'b1101] [18] = 21'h 0007FF;  // +1.9999999999987874 = 2^19 * ln( 1 +  1 * 2^(-19+1) + ( 1^2+-1^2) * 2^(-2*19) )   n = 19   d_n = 1-1i 
assign u[4'b1101] [19] = 21'h 0007FF;  // +1.9999999999996969 = 2^20 * ln( 1 +  1 * 2^(-20+1) + ( 1^2+-1^2) * 2^(-2*20) )   n = 20   d_n = 1-1i 
assign u[4'b1101] [20] = 21'h 0007FF;  // +1.9999999999999243 = 2^21 * ln( 1 +  1 * 2^(-21+1) + ( 1^2+-1^2) * 2^(-2*21) )   n = 21   d_n = 1-1i 
assign u[4'b1101] [21] = 21'h 0007FF;  // +1.9999999999999811 = 2^22 * ln( 1 +  1 * 2^(-22+1) + ( 1^2+-1^2) * 2^(-2*22) )   n = 22   d_n = 1-1i 
assign u[4'b1101] [22] = 21'h 0007FF;  // +1.9999999999999953 = 2^23 * ln( 1 +  1 * 2^(-23+1) + ( 1^2+-1^2) * 2^(-2*23) )   n = 23   d_n = 1-1i 
assign u[4'b1101] [23] = 21'h 0007FF;  // +1.9999999999999989 = 2^24 * ln( 1 +  1 * 2^(-24+1) + ( 1^2+-1^2) * 2^(-2*24) )   n = 24   d_n = 1-1i 
assign u[4'b1101] [24] = 21'h 0007FF;  // +1.9999999999999998 = 2^25 * ln( 1 +  1 * 2^(-25+1) + ( 1^2+-1^2) * 2^(-2*25) )   n = 25   d_n = 1-1i 
assign u[4'b1101] [25] = 21'h 0007FF;  // +1.9999999850988390 = 2^26 * ln( 1 +  1 * 2^(-26+1) + ( 1^2+-1^2) * 2^(-2*26) )   n = 26   d_n = 1-1i 
assign u[4'b1101] [26] = 21'h 0007FF;  // +1.9999999925494194 = 2^27 * ln( 1 +  1 * 2^(-27+1) + ( 1^2+-1^2) * 2^(-2*27) )   n = 27   d_n = 1-1i 
assign u[4'b1101] [27] = 21'h 0007FF;  // +1.9999999962747097 = 2^28 * ln( 1 +  1 * 2^(-28+1) + ( 1^2+-1^2) * 2^(-2*28) )   n = 28   d_n = 1-1i 
assign u[4'b1101] [28] = 21'h 0007FF;  // +1.9999999981373549 = 2^29 * ln( 1 +  1 * 2^(-29+1) + ( 1^2+-1^2) * 2^(-2*29) )   n = 29   d_n = 1-1i 
assign u[4'b1101] [29] = 21'h 0007FF;  // +1.9999999990686774 = 2^30 * ln( 1 +  1 * 2^(-30+1) + ( 1^2+-1^2) * 2^(-2*30) )   n = 30   d_n = 1-1i 
assign u[4'b1101] [30] = 21'h 0007FF;  // +1.9999999995343387 = 2^31 * ln( 1 +  1 * 2^(-31+1) + ( 1^2+-1^2) * 2^(-2*31) )   n = 31   d_n = 1-1i 
assign u[4'b1101] [31] = 21'h 0007FF;  // +1.9999999997671694 = 2^32 * ln( 1 +  1 * 2^(-32+1) + ( 1^2+-1^2) * 2^(-2*32) )   n = 32   d_n = 1-1i 
assign u[4'b1101] [32] = 21'h 0007FF;  // +1.9999999998835847 = 2^33 * ln( 1 +  1 * 2^(-33+1) + ( 1^2+-1^2) * 2^(-2*33) )   n = 33   d_n = 1-1i 
assign u[4'b1101] [33] = 21'h 0007FF;  // +1.9999999999417923 = 2^34 * ln( 1 +  1 * 2^(-34+1) + ( 1^2+-1^2) * 2^(-2*34) )   n = 34   d_n = 1-1i 
assign u[4'b1101] [34] = 21'h 0007FF;  // +1.9999999999708962 = 2^35 * ln( 1 +  1 * 2^(-35+1) + ( 1^2+-1^2) * 2^(-2*35) )   n = 35   d_n = 1-1i 
assign u[4'b1101] [35] = 21'h 0007FF;  // +1.9999999999854481 = 2^36 * ln( 1 +  1 * 2^(-36+1) + ( 1^2+-1^2) * 2^(-2*36) )   n = 36   d_n = 1-1i 
assign u[4'b1101] [36] = 21'h 0007FF;  // +1.9999999999927240 = 2^37 * ln( 1 +  1 * 2^(-37+1) + ( 1^2+-1^2) * 2^(-2*37) )   n = 37   d_n = 1-1i 
assign u[4'b1101] [37] = 21'h 0007FF;  // +1.9999999999963620 = 2^38 * ln( 1 +  1 * 2^(-38+1) + ( 1^2+-1^2) * 2^(-2*38) )   n = 38   d_n = 1-1i 
assign u[4'b1101] [38] = 21'h 0007FF;  // +1.9999999999981810 = 2^39 * ln( 1 +  1 * 2^(-39+1) + ( 1^2+-1^2) * 2^(-2*39) )   n = 39   d_n = 1-1i 
assign u[4'b1101] [39] = 21'h 0007FF;  // +1.9999999999990905 = 2^40 * ln( 1 +  1 * 2^(-40+1) + ( 1^2+-1^2) * 2^(-2*40) )   n = 40   d_n = 1-1i 
assign u[4'b1101] [40] = 21'h 0007FF;  // +1.9999999999995453 = 2^41 * ln( 1 +  1 * 2^(-41+1) + ( 1^2+-1^2) * 2^(-2*41) )   n = 41   d_n = 1-1i 
assign u[4'b1101] [41] = 21'h 0007FF;  // +1.9999999999997726 = 2^42 * ln( 1 +  1 * 2^(-42+1) + ( 1^2+-1^2) * 2^(-2*42) )   n = 42   d_n = 1-1i 
assign u[4'b1101] [42] = 21'h 0007FF;  // +1.9999999999998863 = 2^43 * ln( 1 +  1 * 2^(-43+1) + ( 1^2+-1^2) * 2^(-2*43) )   n = 43   d_n = 1-1i 
assign u[4'b1101] [43] = 21'h 0007FF;  // +1.9999999999999432 = 2^44 * ln( 1 +  1 * 2^(-44+1) + ( 1^2+-1^2) * 2^(-2*44) )   n = 44   d_n = 1-1i 
assign u[4'b1101] [44] = 21'h 0007FF;  // +1.9999999999999716 = 2^45 * ln( 1 +  1 * 2^(-45+1) + ( 1^2+-1^2) * 2^(-2*45) )   n = 45   d_n = 1-1i 
assign u[4'b1101] [45] = 21'h 0007FF;  // +1.9999999999999858 = 2^46 * ln( 1 +  1 * 2^(-46+1) + ( 1^2+-1^2) * 2^(-2*46) )   n = 46   d_n = 1-1i 
assign u[4'b1101] [46] = 21'h 0007FF;  // +1.9999999999999929 = 2^47 * ln( 1 +  1 * 2^(-47+1) + ( 1^2+-1^2) * 2^(-2*47) )   n = 47   d_n = 1-1i 
assign u[4'b1101] [47] = 21'h 0007FF;  // +1.9999999999999964 = 2^48 * ln( 1 +  1 * 2^(-48+1) + ( 1^2+-1^2) * 2^(-2*48) )   n = 48   d_n = 1-1i 
assign u[4'b1101] [48] = 21'h 0007FF;  // +1.9999999999999982 = 2^49 * ln( 1 +  1 * 2^(-49+1) + ( 1^2+-1^2) * 2^(-2*49) )   n = 49   d_n = 1-1i 
assign u[4'b1101] [49] = 21'h 0007FF;  // +1.9999999999999991 = 2^50 * ln( 1 +  1 * 2^(-50+1) + ( 1^2+-1^2) * 2^(-2*50) )   n = 50   d_n = 1-1i 
assign u[4'b1101] [50] = 21'h 0007FF;  // +1.9999999999999996 = 2^51 * ln( 1 +  1 * 2^(-51+1) + ( 1^2+-1^2) * 2^(-2*51) )   n = 51   d_n = 1-1i 
assign u[4'b1101] [51] = 21'h 0007FF;  // +1.9999999999999998 = 2^52 * ln( 1 +  1 * 2^(-52+1) + ( 1^2+-1^2) * 2^(-2*52) )   n = 52   d_n = 1-1i 
assign u[4'b1101] [52] = 21'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  1 * 2^(-53+1) + ( 1^2+-1^2) * 2^(-2*53) )   n = 53   d_n = 1-1i 
assign u[4'b1101] [53] = 21'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  1 * 2^(-54+1) + ( 1^2+-1^2) * 2^(-2*54) )   n = 54   d_n = 1-1i 
assign u[4'b1101] [54] = 21'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  1 * 2^(-55+1) + ( 1^2+-1^2) * 2^(-2*55) )   n = 55   d_n = 1-1i 
assign u[4'b1101] [55] = 21'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  1 * 2^(-56+1) + ( 1^2+-1^2) * 2^(-2*56) )   n = 56   d_n = 1-1i 
assign u[4'b1101] [56] = 21'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  1 * 2^(-57+1) + ( 1^2+-1^2) * 2^(-2*57) )   n = 57   d_n = 1-1i 
assign u[4'b1101] [57] = 21'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  1 * 2^(-58+1) + ( 1^2+-1^2) * 2^(-2*58) )   n = 58   d_n = 1-1i 
assign u[4'b1101] [58] = 21'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  1 * 2^(-59+1) + ( 1^2+-1^2) * 2^(-2*59) )   n = 59   d_n = 1-1i 
assign u[4'b1101] [59] = 21'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  1 * 2^(-60+1) + ( 1^2+-1^2) * 2^(-2*60) )   n = 60   d_n = 1-1i 
assign u[4'b1101] [60] = 21'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  1 * 2^(-61+1) + ( 1^2+-1^2) * 2^(-2*61) )   n = 61   d_n = 1-1i 
assign u[4'b1101] [61] = 21'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  1 * 2^(-62+1) + ( 1^2+-1^2) * 2^(-2*62) )   n = 62   d_n = 1-1i 
assign u[4'b1101] [62] = 21'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  1 * 2^(-63+1) + ( 1^2+-1^2) * 2^(-2*63) )   n = 63   d_n = 1-1i 
assign u[4'b1101] [63] = 21'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  1 * 2^(-64+1) + ( 1^2+-1^2) * 2^(-2*64) )   n = 64   d_n = 1-1i 
assign u[4'b1110] [00] = 21'h 0001C8;  // +0.4462871026284197 = 2^ 1 * ln( 1 +  0 * 2^(- 1+1) + ( 0^2+-1^2) * 2^(-2* 1) )   n =  1   d_n = -0-1i 
assign u[4'b1110] [01] = 21'h 0000F8;  // +0.2424984872657394 = 2^ 2 * ln( 1 +  0 * 2^(- 2+1) + ( 0^2+-1^2) * 2^(-2* 2) )   n =  2   d_n = -0-1i 
assign u[4'b1110] [02] = 21'h 00007F;  // +0.1240334922877210 = 2^ 3 * ln( 1 +  0 * 2^(- 3+1) + ( 0^2+-1^2) * 2^(-2* 3) )   n =  3   d_n = -0-1i 
assign u[4'b1110] [03] = 21'h 00003F;  // +0.0623782466505195 = 2^ 4 * ln( 1 +  0 * 2^(- 4+1) + ( 0^2+-1^2) * 2^(-2* 4) )   n =  4   d_n = -0-1i 
assign u[4'b1110] [04] = 21'h 00001F;  // +0.0312347511377731 = 2^ 5 * ln( 1 +  0 * 2^(- 5+1) + ( 0^2+-1^2) * 2^(-2* 5) )   n =  5   d_n = -0-1i 
assign u[4'b1110] [05] = 21'h 00000F;  // +0.0156230929617406 = 2^ 6 * ln( 1 +  0 * 2^(- 6+1) + ( 0^2+-1^2) * 2^(-2* 6) )   n =  6   d_n = -0-1i 
assign u[4'b1110] [06] = 21'h 000007;  // +0.0078122615911219 = 2^ 7 * ln( 1 +  0 * 2^(- 7+1) + ( 0^2+-1^2) * 2^(-2* 7) )   n =  7   d_n = -0-1i 
assign u[4'b1110] [07] = 21'h 000003;  // +0.0039062201979808 = 2^ 8 * ln( 1 +  0 * 2^(- 8+1) + ( 0^2+-1^2) * 2^(-2* 8) )   n =  8   d_n = -0-1i 
assign u[4'b1110] [08] = 21'h 000001;  // +0.0019531212747156 = 2^ 9 * ln( 1 +  0 * 2^(- 9+1) + ( 0^2+-1^2) * 2^(-2* 9) )   n =  9   d_n = -0-1i 
assign u[4'b1110] [09] = 21'h 000000;  // +0.0009765620343389 = 2^10 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+-1^2) * 2^(-2*10) )   n = 10   d_n = -0-1i 
assign u[4'b1110] [10] = 21'h 000000;  // +0.0004882811917923 = 2^11 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+-1^2) * 2^(-2*11) )   n = 11   d_n = -0-1i 
assign u[4'b1110] [11] = 21'h 000000;  // +0.0002441406177240 = 2^12 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+-1^2) * 2^(-2*12) )   n = 12   d_n = -0-1i 
assign u[4'b1110] [12] = 21'h 000000;  // +0.0001220703120453 = 2^13 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+-1^2) * 2^(-2*13) )   n = 13   d_n = -0-1i 
assign u[4'b1110] [13] = 21'h 000000;  // +0.0000610351561932 = 2^14 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+-1^2) * 2^(-2*14) )   n = 14   d_n = -0-1i 
assign u[4'b1110] [14] = 21'h 000000;  // +0.0000305175781179 = 2^15 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+-1^2) * 2^(-2*15) )   n = 15   d_n = -0-1i 
assign u[4'b1110] [15] = 21'h 000000;  // +0.0000152587890616 = 2^16 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+-1^2) * 2^(-2*16) )   n = 16   d_n = -0-1i 
assign u[4'b1110] [16] = 21'h 000000;  // +0.0000076293945311 = 2^17 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+-1^2) * 2^(-2*17) )   n = 17   d_n = -0-1i 
assign u[4'b1110] [17] = 21'h 000000;  // +0.0000038146972656 = 2^18 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+-1^2) * 2^(-2*18) )   n = 18   d_n = -0-1i 
assign u[4'b1110] [18] = 21'h 000000;  // +0.0000019073486328 = 2^19 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+-1^2) * 2^(-2*19) )   n = 19   d_n = -0-1i 
assign u[4'b1110] [19] = 21'h 000000;  // +0.0000009536743164 = 2^20 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+-1^2) * 2^(-2*20) )   n = 20   d_n = -0-1i 
assign u[4'b1110] [20] = 21'h 000000;  // +0.0000004768371582 = 2^21 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+-1^2) * 2^(-2*21) )   n = 21   d_n = -0-1i 
assign u[4'b1110] [21] = 21'h 000000;  // +0.0000002384185791 = 2^22 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+-1^2) * 2^(-2*22) )   n = 22   d_n = -0-1i 
assign u[4'b1110] [22] = 21'h 000000;  // +0.0000001192092896 = 2^23 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+-1^2) * 2^(-2*23) )   n = 23   d_n = -0-1i 
assign u[4'b1110] [23] = 21'h 000000;  // +0.0000000596046448 = 2^24 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+-1^2) * 2^(-2*24) )   n = 24   d_n = -0-1i 
assign u[4'b1110] [24] = 21'h 000000;  // +0.0000000298023224 = 2^25 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+-1^2) * 2^(-2*25) )   n = 25   d_n = -0-1i 
assign u[4'b1110] [25] = 21'h 000000;  // +0.0000000000000000 = 2^26 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+-1^2) * 2^(-2*26) )   n = 26   d_n = -0-1i 
assign u[4'b1110] [26] = 21'h 000000;  // +0.0000000000000000 = 2^27 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+-1^2) * 2^(-2*27) )   n = 27   d_n = -0-1i 
assign u[4'b1110] [27] = 21'h 000000;  // +0.0000000000000000 = 2^28 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+-1^2) * 2^(-2*28) )   n = 28   d_n = -0-1i 
assign u[4'b1110] [28] = 21'h 000000;  // +0.0000000000000000 = 2^29 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+-1^2) * 2^(-2*29) )   n = 29   d_n = -0-1i 
assign u[4'b1110] [29] = 21'h 000000;  // +0.0000000000000000 = 2^30 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+-1^2) * 2^(-2*30) )   n = 30   d_n = -0-1i 
assign u[4'b1110] [30] = 21'h 000000;  // +0.0000000000000000 = 2^31 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+-1^2) * 2^(-2*31) )   n = 31   d_n = -0-1i 
assign u[4'b1110] [31] = 21'h 000000;  // +0.0000000000000000 = 2^32 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+-1^2) * 2^(-2*32) )   n = 32   d_n = -0-1i 
assign u[4'b1110] [32] = 21'h 000000;  // +0.0000000000000000 = 2^33 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+-1^2) * 2^(-2*33) )   n = 33   d_n = -0-1i 
assign u[4'b1110] [33] = 21'h 000000;  // +0.0000000000000000 = 2^34 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+-1^2) * 2^(-2*34) )   n = 34   d_n = -0-1i 
assign u[4'b1110] [34] = 21'h 000000;  // +0.0000000000000000 = 2^35 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+-1^2) * 2^(-2*35) )   n = 35   d_n = -0-1i 
assign u[4'b1110] [35] = 21'h 000000;  // +0.0000000000000000 = 2^36 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+-1^2) * 2^(-2*36) )   n = 36   d_n = -0-1i 
assign u[4'b1110] [36] = 21'h 000000;  // +0.0000000000000000 = 2^37 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+-1^2) * 2^(-2*37) )   n = 37   d_n = -0-1i 
assign u[4'b1110] [37] = 21'h 000000;  // +0.0000000000000000 = 2^38 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+-1^2) * 2^(-2*38) )   n = 38   d_n = -0-1i 
assign u[4'b1110] [38] = 21'h 000000;  // +0.0000000000000000 = 2^39 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+-1^2) * 2^(-2*39) )   n = 39   d_n = -0-1i 
assign u[4'b1110] [39] = 21'h 000000;  // +0.0000000000000000 = 2^40 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+-1^2) * 2^(-2*40) )   n = 40   d_n = -0-1i 
assign u[4'b1110] [40] = 21'h 000000;  // +0.0000000000000000 = 2^41 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+-1^2) * 2^(-2*41) )   n = 41   d_n = -0-1i 
assign u[4'b1110] [41] = 21'h 000000;  // +0.0000000000000000 = 2^42 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+-1^2) * 2^(-2*42) )   n = 42   d_n = -0-1i 
assign u[4'b1110] [42] = 21'h 000000;  // +0.0000000000000000 = 2^43 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+-1^2) * 2^(-2*43) )   n = 43   d_n = -0-1i 
assign u[4'b1110] [43] = 21'h 000000;  // +0.0000000000000000 = 2^44 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+-1^2) * 2^(-2*44) )   n = 44   d_n = -0-1i 
assign u[4'b1110] [44] = 21'h 000000;  // +0.0000000000000000 = 2^45 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+-1^2) * 2^(-2*45) )   n = 45   d_n = -0-1i 
assign u[4'b1110] [45] = 21'h 000000;  // +0.0000000000000000 = 2^46 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+-1^2) * 2^(-2*46) )   n = 46   d_n = -0-1i 
assign u[4'b1110] [46] = 21'h 000000;  // +0.0000000000000000 = 2^47 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+-1^2) * 2^(-2*47) )   n = 47   d_n = -0-1i 
assign u[4'b1110] [47] = 21'h 000000;  // +0.0000000000000000 = 2^48 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+-1^2) * 2^(-2*48) )   n = 48   d_n = -0-1i 
assign u[4'b1110] [48] = 21'h 000000;  // +0.0000000000000000 = 2^49 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+-1^2) * 2^(-2*49) )   n = 49   d_n = -0-1i 
assign u[4'b1110] [49] = 21'h 000000;  // +0.0000000000000000 = 2^50 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+-1^2) * 2^(-2*50) )   n = 50   d_n = -0-1i 
assign u[4'b1110] [50] = 21'h 000000;  // +0.0000000000000000 = 2^51 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+-1^2) * 2^(-2*51) )   n = 51   d_n = -0-1i 
assign u[4'b1110] [51] = 21'h 000000;  // +0.0000000000000000 = 2^52 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+-1^2) * 2^(-2*52) )   n = 52   d_n = -0-1i 
assign u[4'b1110] [52] = 21'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+-1^2) * 2^(-2*53) )   n = 53   d_n = -0-1i 
assign u[4'b1110] [53] = 21'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+-1^2) * 2^(-2*54) )   n = 54   d_n = -0-1i 
assign u[4'b1110] [54] = 21'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+-1^2) * 2^(-2*55) )   n = 55   d_n = -0-1i 
assign u[4'b1110] [55] = 21'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+-1^2) * 2^(-2*56) )   n = 56   d_n = -0-1i 
assign u[4'b1110] [56] = 21'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+-1^2) * 2^(-2*57) )   n = 57   d_n = -0-1i 
assign u[4'b1110] [57] = 21'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+-1^2) * 2^(-2*58) )   n = 58   d_n = -0-1i 
assign u[4'b1110] [58] = 21'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+-1^2) * 2^(-2*59) )   n = 59   d_n = -0-1i 
assign u[4'b1110] [59] = 21'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+-1^2) * 2^(-2*60) )   n = 60   d_n = -0-1i 
assign u[4'b1110] [60] = 21'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+-1^2) * 2^(-2*61) )   n = 61   d_n = -0-1i 
assign u[4'b1110] [61] = 21'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+-1^2) * 2^(-2*62) )   n = 62   d_n = -0-1i 
assign u[4'b1110] [62] = 21'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+-1^2) * 2^(-2*63) )   n = 63   d_n = -0-1i 
assign u[4'b1110] [63] = 21'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+-1^2) * 2^(-2*64) )   n = 64   d_n = -0-1i 
assign u[4'b1111] [00] = 21'h 1FFA74;  // -1.3862943611198904 = 2^ 1 * ln( 1 + -1 * 2^(- 1+1) + (-1^2+-1^2) * 2^(-2* 1) )   n =  1   d_n = -1-1i 
assign u[4'b1111] [01] = 21'h 1FF87A;  // -1.8800145169829416 = 2^ 2 * ln( 1 + -1 * 2^(- 2+1) + (-1^2+-1^2) * 2^(-2* 2) )   n =  2   d_n = -1-1i 
assign u[4'b1111] [02] = 21'h 1FF819;  // -1.9748806234522058 = 2^ 3 * ln( 1 + -1 * 2^(- 3+1) + (-1^2+-1^2) * 2^(-2* 3) )   n =  3   d_n = -1-1i 
assign u[4'b1111] [03] = 21'h 1FF805;  // -1.9942791233164259 = 2^ 4 * ln( 1 + -1 * 2^(- 4+1) + (-1^2+-1^2) * 2^(-2* 4) )   n =  4   d_n = -1-1i 
assign u[4'b1111] [04] = 21'h 1FF801;  // -1.9986353578798890 = 2^ 5 * ln( 1 + -1 * 2^(- 5+1) + (-1^2+-1^2) * 2^(-2* 5) )   n =  5   d_n = -1-1i 
assign u[4'b1111] [05] = 21'h 1FF800;  // -1.9996667544388824 = 2^ 6 * ln( 1 + -1 * 2^(- 6+1) + (-1^2+-1^2) * 2^(-2* 6) )   n =  6   d_n = -1-1i 
assign u[4'b1111] [06] = 21'h 1FF800;  // -1.9999176601574109 = 2^ 7 * ln( 1 + -1 * 2^(- 7+1) + (-1^2+-1^2) * 2^(-2* 7) )   n =  7   d_n = -1-1i 
assign u[4'b1111] [07] = 21'h 1FF800;  // -1.9999795353661032 = 2^ 8 * ln( 1 + -1 * 2^(- 8+1) + (-1^2+-1^2) * 2^(-2* 8) )   n =  8   d_n = -1-1i 
assign u[4'b1111] [08] = 21'h 1FF800;  // -1.9999948988125242 = 2^ 9 * ln( 1 + -1 * 2^(- 9+1) + (-1^2+-1^2) * 2^(-2* 9) )   n =  9   d_n = -1-1i 
assign u[4'b1111] [09] = 21'h 1FF800;  // -1.9999987265701442 = 2^10 * ln( 1 + -1 * 2^(-10+1) + (-1^2+-1^2) * 2^(-2*10) )   n = 10   d_n = -1-1i 
assign u[4'b1111] [10] = 21'h 1FF800;  // -1.9999996818756538 = 2^11 * ln( 1 + -1 * 2^(-11+1) + (-1^2+-1^2) * 2^(-2*11) )   n = 11   d_n = -1-1i 
assign u[4'b1111] [11] = 21'h 1FF800;  // -1.9999999204980317 = 2^12 * ln( 1 + -1 * 2^(-12+1) + (-1^2+-1^2) * 2^(-2*12) )   n = 12   d_n = -1-1i 
assign u[4'b1111] [12] = 21'h 1FF800;  // -1.9999999801276920 = 2^13 * ln( 1 + -1 * 2^(-13+1) + (-1^2+-1^2) * 2^(-2*13) )   n = 13   d_n = -1-1i 
assign u[4'b1111] [13] = 21'h 1FF800;  // -1.9999999950326621 = 2^14 * ln( 1 + -1 * 2^(-14+1) + (-1^2+-1^2) * 2^(-2*14) )   n = 14   d_n = -1-1i 
assign u[4'b1111] [14] = 21'h 1FF800;  // -1.9999999987582011 = 2^15 * ln( 1 + -1 * 2^(-15+1) + (-1^2+-1^2) * 2^(-2*15) )   n = 15   d_n = -1-1i 
assign u[4'b1111] [15] = 21'h 1FF800;  // -1.9999999996895548 = 2^16 * ln( 1 + -1 * 2^(-16+1) + (-1^2+-1^2) * 2^(-2*16) )   n = 16   d_n = -1-1i 
assign u[4'b1111] [16] = 21'h 1FF800;  // -1.9999999999223892 = 2^17 * ln( 1 + -1 * 2^(-17+1) + (-1^2+-1^2) * 2^(-2*17) )   n = 17   d_n = -1-1i 
assign u[4'b1111] [17] = 21'h 1FF800;  // -1.9999999999951494 = 2^18 * ln( 1 + -1 * 2^(-18+1) + (-1^2+-1^2) * 2^(-2*18) )   n = 18   d_n = -1-1i 
assign u[4'b1111] [18] = 21'h 1FF800;  // -1.9999999999987874 = 2^19 * ln( 1 + -1 * 2^(-19+1) + (-1^2+-1^2) * 2^(-2*19) )   n = 19   d_n = -1-1i 
assign u[4'b1111] [19] = 21'h 1FF800;  // -1.9999999999996969 = 2^20 * ln( 1 + -1 * 2^(-20+1) + (-1^2+-1^2) * 2^(-2*20) )   n = 20   d_n = -1-1i 
assign u[4'b1111] [20] = 21'h 1FF800;  // -1.9999999999999243 = 2^21 * ln( 1 + -1 * 2^(-21+1) + (-1^2+-1^2) * 2^(-2*21) )   n = 21   d_n = -1-1i 
assign u[4'b1111] [21] = 21'h 1FF800;  // -1.9999999999999811 = 2^22 * ln( 1 + -1 * 2^(-22+1) + (-1^2+-1^2) * 2^(-2*22) )   n = 22   d_n = -1-1i 
assign u[4'b1111] [22] = 21'h 1FF800;  // -1.9999999999999953 = 2^23 * ln( 1 + -1 * 2^(-23+1) + (-1^2+-1^2) * 2^(-2*23) )   n = 23   d_n = -1-1i 
assign u[4'b1111] [23] = 21'h 1FF800;  // -1.9999999999999989 = 2^24 * ln( 1 + -1 * 2^(-24+1) + (-1^2+-1^2) * 2^(-2*24) )   n = 24   d_n = -1-1i 
assign u[4'b1111] [24] = 21'h 1FF800;  // -1.9999999999999998 = 2^25 * ln( 1 + -1 * 2^(-25+1) + (-1^2+-1^2) * 2^(-2*25) )   n = 25   d_n = -1-1i 
assign u[4'b1111] [25] = 21'h 1FF800;  // -2.0000000000000000 = 2^26 * ln( 1 + -1 * 2^(-26+1) + (-1^2+-1^2) * 2^(-2*26) )   n = 26   d_n = -1-1i 
assign u[4'b1111] [26] = 21'h 1FF7FF;  // -2.0000000074505806 = 2^27 * ln( 1 + -1 * 2^(-27+1) + (-1^2+-1^2) * 2^(-2*27) )   n = 27   d_n = -1-1i 
assign u[4'b1111] [27] = 21'h 1FF7FF;  // -2.0000000037252903 = 2^28 * ln( 1 + -1 * 2^(-28+1) + (-1^2+-1^2) * 2^(-2*28) )   n = 28   d_n = -1-1i 
assign u[4'b1111] [28] = 21'h 1FF7FF;  // -2.0000000018626451 = 2^29 * ln( 1 + -1 * 2^(-29+1) + (-1^2+-1^2) * 2^(-2*29) )   n = 29   d_n = -1-1i 
assign u[4'b1111] [29] = 21'h 1FF7FF;  // -2.0000000009313226 = 2^30 * ln( 1 + -1 * 2^(-30+1) + (-1^2+-1^2) * 2^(-2*30) )   n = 30   d_n = -1-1i 
assign u[4'b1111] [30] = 21'h 1FF7FF;  // -2.0000000004656613 = 2^31 * ln( 1 + -1 * 2^(-31+1) + (-1^2+-1^2) * 2^(-2*31) )   n = 31   d_n = -1-1i 
assign u[4'b1111] [31] = 21'h 1FF7FF;  // -2.0000000002328306 = 2^32 * ln( 1 + -1 * 2^(-32+1) + (-1^2+-1^2) * 2^(-2*32) )   n = 32   d_n = -1-1i 
assign u[4'b1111] [32] = 21'h 1FF7FF;  // -2.0000000001164153 = 2^33 * ln( 1 + -1 * 2^(-33+1) + (-1^2+-1^2) * 2^(-2*33) )   n = 33   d_n = -1-1i 
assign u[4'b1111] [33] = 21'h 1FF7FF;  // -2.0000000000582077 = 2^34 * ln( 1 + -1 * 2^(-34+1) + (-1^2+-1^2) * 2^(-2*34) )   n = 34   d_n = -1-1i 
assign u[4'b1111] [34] = 21'h 1FF7FF;  // -2.0000000000291038 = 2^35 * ln( 1 + -1 * 2^(-35+1) + (-1^2+-1^2) * 2^(-2*35) )   n = 35   d_n = -1-1i 
assign u[4'b1111] [35] = 21'h 1FF7FF;  // -2.0000000000145519 = 2^36 * ln( 1 + -1 * 2^(-36+1) + (-1^2+-1^2) * 2^(-2*36) )   n = 36   d_n = -1-1i 
assign u[4'b1111] [36] = 21'h 1FF7FF;  // -2.0000000000072760 = 2^37 * ln( 1 + -1 * 2^(-37+1) + (-1^2+-1^2) * 2^(-2*37) )   n = 37   d_n = -1-1i 
assign u[4'b1111] [37] = 21'h 1FF7FF;  // -2.0000000000036380 = 2^38 * ln( 1 + -1 * 2^(-38+1) + (-1^2+-1^2) * 2^(-2*38) )   n = 38   d_n = -1-1i 
assign u[4'b1111] [38] = 21'h 1FF7FF;  // -2.0000000000018190 = 2^39 * ln( 1 + -1 * 2^(-39+1) + (-1^2+-1^2) * 2^(-2*39) )   n = 39   d_n = -1-1i 
assign u[4'b1111] [39] = 21'h 1FF7FF;  // -2.0000000000009095 = 2^40 * ln( 1 + -1 * 2^(-40+1) + (-1^2+-1^2) * 2^(-2*40) )   n = 40   d_n = -1-1i 
assign u[4'b1111] [40] = 21'h 1FF7FF;  // -2.0000000000004547 = 2^41 * ln( 1 + -1 * 2^(-41+1) + (-1^2+-1^2) * 2^(-2*41) )   n = 41   d_n = -1-1i 
assign u[4'b1111] [41] = 21'h 1FF7FF;  // -2.0000000000002274 = 2^42 * ln( 1 + -1 * 2^(-42+1) + (-1^2+-1^2) * 2^(-2*42) )   n = 42   d_n = -1-1i 
assign u[4'b1111] [42] = 21'h 1FF800;  // -2.0000000000001137 = 2^43 * ln( 1 + -1 * 2^(-43+1) + (-1^2+-1^2) * 2^(-2*43) )   n = 43   d_n = -1-1i 
assign u[4'b1111] [43] = 21'h 1FF800;  // -2.0000000000000568 = 2^44 * ln( 1 + -1 * 2^(-44+1) + (-1^2+-1^2) * 2^(-2*44) )   n = 44   d_n = -1-1i 
assign u[4'b1111] [44] = 21'h 1FF800;  // -2.0000000000000284 = 2^45 * ln( 1 + -1 * 2^(-45+1) + (-1^2+-1^2) * 2^(-2*45) )   n = 45   d_n = -1-1i 
assign u[4'b1111] [45] = 21'h 1FF800;  // -2.0000000000000142 = 2^46 * ln( 1 + -1 * 2^(-46+1) + (-1^2+-1^2) * 2^(-2*46) )   n = 46   d_n = -1-1i 
assign u[4'b1111] [46] = 21'h 1FF800;  // -2.0000000000000071 = 2^47 * ln( 1 + -1 * 2^(-47+1) + (-1^2+-1^2) * 2^(-2*47) )   n = 47   d_n = -1-1i 
assign u[4'b1111] [47] = 21'h 1FF800;  // -2.0000000000000036 = 2^48 * ln( 1 + -1 * 2^(-48+1) + (-1^2+-1^2) * 2^(-2*48) )   n = 48   d_n = -1-1i 
assign u[4'b1111] [48] = 21'h 1FF800;  // -2.0000000000000018 = 2^49 * ln( 1 + -1 * 2^(-49+1) + (-1^2+-1^2) * 2^(-2*49) )   n = 49   d_n = -1-1i 
assign u[4'b1111] [49] = 21'h 1FF800;  // -2.0000000000000009 = 2^50 * ln( 1 + -1 * 2^(-50+1) + (-1^2+-1^2) * 2^(-2*50) )   n = 50   d_n = -1-1i 
assign u[4'b1111] [50] = 21'h 1FF800;  // -2.0000000000000004 = 2^51 * ln( 1 + -1 * 2^(-51+1) + (-1^2+-1^2) * 2^(-2*51) )   n = 51   d_n = -1-1i 
assign u[4'b1111] [51] = 21'h 1FF800;  // -2.0000000000000004 = 2^52 * ln( 1 + -1 * 2^(-52+1) + (-1^2+-1^2) * 2^(-2*52) )   n = 52   d_n = -1-1i 
assign u[4'b1111] [52] = 21'h 1FF800;  // -2.0000000000000000 = 2^53 * ln( 1 + -1 * 2^(-53+1) + (-1^2+-1^2) * 2^(-2*53) )   n = 53   d_n = -1-1i 
assign u[4'b1111] [53] = 21'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 + -1 * 2^(-54+1) + (-1^2+-1^2) * 2^(-2*54) )   n = 54   d_n = -1-1i 
assign u[4'b1111] [54] = 21'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 + -1 * 2^(-55+1) + (-1^2+-1^2) * 2^(-2*55) )   n = 55   d_n = -1-1i 
assign u[4'b1111] [55] = 21'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 + -1 * 2^(-56+1) + (-1^2+-1^2) * 2^(-2*56) )   n = 56   d_n = -1-1i 
assign u[4'b1111] [56] = 21'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 + -1 * 2^(-57+1) + (-1^2+-1^2) * 2^(-2*57) )   n = 57   d_n = -1-1i 
assign u[4'b1111] [57] = 21'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 + -1 * 2^(-58+1) + (-1^2+-1^2) * 2^(-2*58) )   n = 58   d_n = -1-1i 
assign u[4'b1111] [58] = 21'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 + -1 * 2^(-59+1) + (-1^2+-1^2) * 2^(-2*59) )   n = 59   d_n = -1-1i 
assign u[4'b1111] [59] = 21'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 + -1 * 2^(-60+1) + (-1^2+-1^2) * 2^(-2*60) )   n = 60   d_n = -1-1i 
assign u[4'b1111] [60] = 21'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 + -1 * 2^(-61+1) + (-1^2+-1^2) * 2^(-2*61) )   n = 61   d_n = -1-1i 
assign u[4'b1111] [61] = 21'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 + -1 * 2^(-62+1) + (-1^2+-1^2) * 2^(-2*62) )   n = 62   d_n = -1-1i 
assign u[4'b1111] [62] = 21'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 + -1 * 2^(-63+1) + (-1^2+-1^2) * 2^(-2*63) )   n = 63   d_n = -1-1i 
assign u[4'b1111] [63] = 21'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 + -1 * 2^(-64+1) + (-1^2+-1^2) * 2^(-2*64) )   n = 64   d_n = -1-1i 
assign v[4'b0000] [00] = 21'h 000000;  // +0.0000000000000000 = 2^(1+1) *  0 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = 0 
assign v[4'b0000] [01] = 21'h 000000;  // +0.0000000000000000 = 2^(2+1) *  0 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = 0 
assign v[4'b0000] [02] = 21'h 000000;  // +0.0000000000000000 = 2^(3+1) *  0 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = 0 
assign v[4'b0000] [03] = 21'h 000000;  // +0.0000000000000000 = 2^(4+1) *  0 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = 0 
assign v[4'b0000] [04] = 21'h 000000;  // +0.0000000000000000 = 2^(5+1) *  0 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = 0 
assign v[4'b0000] [05] = 21'h 000000;  // +0.0000000000000000 = 2^(6+1) *  0 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = 0 
assign v[4'b0000] [06] = 21'h 000000;  // +0.0000000000000000 = 2^(7+1) *  0 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = 0 
assign v[4'b0000] [07] = 21'h 000000;  // +0.0000000000000000 = 2^(8+1) *  0 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = 0 
assign v[4'b0000] [08] = 21'h 000000;  // +0.0000000000000000 = 2^(9+1) *  0 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = 0 
assign v[4'b0000] [09] = 21'h 000000;  // +0.0000000000000000 = 2^(10+1) *  0 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = 0 
assign v[4'b0000] [10] = 21'h 000000;  // +0.0000000000000000 = 2^(11+1) *  0 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = 0 
assign v[4'b0000] [11] = 21'h 000000;  // +0.0000000000000000 = 2^(12+1) *  0 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = 0 
assign v[4'b0000] [12] = 21'h 000000;  // +0.0000000000000000 = 2^(13+1) *  0 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = 0 
assign v[4'b0000] [13] = 21'h 000000;  // +0.0000000000000000 = 2^(14+1) *  0 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = 0 
assign v[4'b0000] [14] = 21'h 000000;  // +0.0000000000000000 = 2^(15+1) *  0 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = 0 
assign v[4'b0000] [15] = 21'h 000000;  // +0.0000000000000000 = 2^(16+1) *  0 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = 0 
assign v[4'b0000] [16] = 21'h 000000;  // +0.0000000000000000 = 2^(17+1) *  0 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = 0 
assign v[4'b0000] [17] = 21'h 000000;  // +0.0000000000000000 = 2^(18+1) *  0 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = 0 
assign v[4'b0000] [18] = 21'h 000000;  // +0.0000000000000000 = 2^(19+1) *  0 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = 0 
assign v[4'b0000] [19] = 21'h 000000;  // +0.0000000000000000 = 2^(20+1) *  0 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = 0 
assign v[4'b0000] [20] = 21'h 000000;  // +0.0000000000000000 = 2^(21+1) *  0 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = 0 
assign v[4'b0000] [21] = 21'h 000000;  // +0.0000000000000000 = 2^(22+1) *  0 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = 0 
assign v[4'b0000] [22] = 21'h 000000;  // +0.0000000000000000 = 2^(23+1) *  0 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = 0 
assign v[4'b0000] [23] = 21'h 000000;  // +0.0000000000000000 = 2^(24+1) *  0 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = 0 
assign v[4'b0000] [24] = 21'h 000000;  // +0.0000000000000000 = 2^(25+1) *  0 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = 0 
assign v[4'b0000] [25] = 21'h 000000;  // +0.0000000000000000 = 2^(26+1) *  0 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = 0 
assign v[4'b0000] [26] = 21'h 000000;  // +0.0000000000000000 = 2^(27+1) *  0 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = 0 
assign v[4'b0000] [27] = 21'h 000000;  // +0.0000000000000000 = 2^(28+1) *  0 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = 0 
assign v[4'b0000] [28] = 21'h 000000;  // +0.0000000000000000 = 2^(29+1) *  0 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = 0 
assign v[4'b0000] [29] = 21'h 000000;  // +0.0000000000000000 = 2^(30+1) *  0 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = 0 
assign v[4'b0000] [30] = 21'h 000000;  // +0.0000000000000000 = 2^(31+1) *  0 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = 0 
assign v[4'b0000] [31] = 21'h 000000;  // +0.0000000000000000 = 2^(32+1) *  0 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = 0 
assign v[4'b0000] [32] = 21'h 000000;  // +0.0000000000000000 = 2^(33+1) *  0 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = 0 
assign v[4'b0000] [33] = 21'h 000000;  // +0.0000000000000000 = 2^(34+1) *  0 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = 0 
assign v[4'b0000] [34] = 21'h 000000;  // +0.0000000000000000 = 2^(35+1) *  0 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = 0 
assign v[4'b0000] [35] = 21'h 000000;  // +0.0000000000000000 = 2^(36+1) *  0 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = 0 
assign v[4'b0000] [36] = 21'h 000000;  // +0.0000000000000000 = 2^(37+1) *  0 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = 0 
assign v[4'b0000] [37] = 21'h 000000;  // +0.0000000000000000 = 2^(38+1) *  0 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = 0 
assign v[4'b0000] [38] = 21'h 000000;  // +0.0000000000000000 = 2^(39+1) *  0 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = 0 
assign v[4'b0000] [39] = 21'h 000000;  // +0.0000000000000000 = 2^(40+1) *  0 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = 0 
assign v[4'b0000] [40] = 21'h 000000;  // +0.0000000000000000 = 2^(41+1) *  0 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = 0 
assign v[4'b0000] [41] = 21'h 000000;  // +0.0000000000000000 = 2^(42+1) *  0 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = 0 
assign v[4'b0000] [42] = 21'h 000000;  // +0.0000000000000000 = 2^(43+1) *  0 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = 0 
assign v[4'b0000] [43] = 21'h 000000;  // +0.0000000000000000 = 2^(44+1) *  0 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = 0 
assign v[4'b0000] [44] = 21'h 000000;  // +0.0000000000000000 = 2^(45+1) *  0 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = 0 
assign v[4'b0000] [45] = 21'h 000000;  // +0.0000000000000000 = 2^(46+1) *  0 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = 0 
assign v[4'b0000] [46] = 21'h 000000;  // +0.0000000000000000 = 2^(47+1) *  0 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = 0 
assign v[4'b0000] [47] = 21'h 000000;  // +0.0000000000000000 = 2^(48+1) *  0 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = 0 
assign v[4'b0000] [48] = 21'h 000000;  // +0.0000000000000000 = 2^(49+1) *  0 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = 0 
assign v[4'b0000] [49] = 21'h 000000;  // +0.0000000000000000 = 2^(50+1) *  0 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = 0 
assign v[4'b0000] [50] = 21'h 000000;  // +0.0000000000000000 = 2^(51+1) *  0 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = 0 
assign v[4'b0000] [51] = 21'h 000000;  // +0.0000000000000000 = 2^(52+1) *  0 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = 0 
assign v[4'b0000] [52] = 21'h 000000;  // +0.0000000000000000 = 2^(53+1) *  0 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = 0 
assign v[4'b0000] [53] = 21'h 000000;  // +0.0000000000000000 = 2^(54+1) *  0 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = 0 
assign v[4'b0000] [54] = 21'h 000000;  // +0.0000000000000000 = 2^(55+1) *  0 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = 0 
assign v[4'b0000] [55] = 21'h 000000;  // +0.0000000000000000 = 2^(56+1) *  0 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = 0 
assign v[4'b0000] [56] = 21'h 000000;  // +0.0000000000000000 = 2^(57+1) *  0 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = 0 
assign v[4'b0000] [57] = 21'h 000000;  // +0.0000000000000000 = 2^(58+1) *  0 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = 0 
assign v[4'b0000] [58] = 21'h 000000;  // +0.0000000000000000 = 2^(59+1) *  0 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = 0 
assign v[4'b0000] [59] = 21'h 000000;  // +0.0000000000000000 = 2^(60+1) *  0 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = 0 
assign v[4'b0000] [60] = 21'h 000000;  // +0.0000000000000000 = 2^(61+1) *  0 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = 0 
assign v[4'b0000] [61] = 21'h 000000;  // +0.0000000000000000 = 2^(62+1) *  0 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = 0 
assign v[4'b0000] [62] = 21'h 000000;  // +0.0000000000000000 = 2^(63+1) *  0 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = 0 
assign v[4'b0000] [63] = 21'h 000000;  // +0.0000000000000000 = 2^(64+1) *  0 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = 0 
assign v[4'b0001] [00] = 21'h 000000;  // +0.0000000000000000 = 2^(1+1) *  0 * atan( 1 / (  1 + 2^1 ) )   n =  1   d_n = 1 
assign v[4'b0001] [01] = 21'h 000000;  // +0.0000000000000000 = 2^(2+1) *  0 * atan( 1 / (  1 + 2^2 ) )   n =  2   d_n = 1 
assign v[4'b0001] [02] = 21'h 000000;  // +0.0000000000000000 = 2^(3+1) *  0 * atan( 1 / (  1 + 2^3 ) )   n =  3   d_n = 1 
assign v[4'b0001] [03] = 21'h 000000;  // +0.0000000000000000 = 2^(4+1) *  0 * atan( 1 / (  1 + 2^4 ) )   n =  4   d_n = 1 
assign v[4'b0001] [04] = 21'h 000000;  // +0.0000000000000000 = 2^(5+1) *  0 * atan( 1 / (  1 + 2^5 ) )   n =  5   d_n = 1 
assign v[4'b0001] [05] = 21'h 000000;  // +0.0000000000000000 = 2^(6+1) *  0 * atan( 1 / (  1 + 2^6 ) )   n =  6   d_n = 1 
assign v[4'b0001] [06] = 21'h 000000;  // +0.0000000000000000 = 2^(7+1) *  0 * atan( 1 / (  1 + 2^7 ) )   n =  7   d_n = 1 
assign v[4'b0001] [07] = 21'h 000000;  // +0.0000000000000000 = 2^(8+1) *  0 * atan( 1 / (  1 + 2^8 ) )   n =  8   d_n = 1 
assign v[4'b0001] [08] = 21'h 000000;  // +0.0000000000000000 = 2^(9+1) *  0 * atan( 1 / (  1 + 2^9 ) )   n =  9   d_n = 1 
assign v[4'b0001] [09] = 21'h 000000;  // +0.0000000000000000 = 2^(10+1) *  0 * atan( 1 / (  1 + 2^10 ) )   n = 10   d_n = 1 
assign v[4'b0001] [10] = 21'h 000000;  // +0.0000000000000000 = 2^(11+1) *  0 * atan( 1 / (  1 + 2^11 ) )   n = 11   d_n = 1 
assign v[4'b0001] [11] = 21'h 000000;  // +0.0000000000000000 = 2^(12+1) *  0 * atan( 1 / (  1 + 2^12 ) )   n = 12   d_n = 1 
assign v[4'b0001] [12] = 21'h 000000;  // +0.0000000000000000 = 2^(13+1) *  0 * atan( 1 / (  1 + 2^13 ) )   n = 13   d_n = 1 
assign v[4'b0001] [13] = 21'h 000000;  // +0.0000000000000000 = 2^(14+1) *  0 * atan( 1 / (  1 + 2^14 ) )   n = 14   d_n = 1 
assign v[4'b0001] [14] = 21'h 000000;  // +0.0000000000000000 = 2^(15+1) *  0 * atan( 1 / (  1 + 2^15 ) )   n = 15   d_n = 1 
assign v[4'b0001] [15] = 21'h 000000;  // +0.0000000000000000 = 2^(16+1) *  0 * atan( 1 / (  1 + 2^16 ) )   n = 16   d_n = 1 
assign v[4'b0001] [16] = 21'h 000000;  // +0.0000000000000000 = 2^(17+1) *  0 * atan( 1 / (  1 + 2^17 ) )   n = 17   d_n = 1 
assign v[4'b0001] [17] = 21'h 000000;  // +0.0000000000000000 = 2^(18+1) *  0 * atan( 1 / (  1 + 2^18 ) )   n = 18   d_n = 1 
assign v[4'b0001] [18] = 21'h 000000;  // +0.0000000000000000 = 2^(19+1) *  0 * atan( 1 / (  1 + 2^19 ) )   n = 19   d_n = 1 
assign v[4'b0001] [19] = 21'h 000000;  // +0.0000000000000000 = 2^(20+1) *  0 * atan( 1 / (  1 + 2^20 ) )   n = 20   d_n = 1 
assign v[4'b0001] [20] = 21'h 000000;  // +0.0000000000000000 = 2^(21+1) *  0 * atan( 1 / (  1 + 2^21 ) )   n = 21   d_n = 1 
assign v[4'b0001] [21] = 21'h 000000;  // +0.0000000000000000 = 2^(22+1) *  0 * atan( 1 / (  1 + 2^22 ) )   n = 22   d_n = 1 
assign v[4'b0001] [22] = 21'h 000000;  // +0.0000000000000000 = 2^(23+1) *  0 * atan( 1 / (  1 + 2^23 ) )   n = 23   d_n = 1 
assign v[4'b0001] [23] = 21'h 000000;  // +0.0000000000000000 = 2^(24+1) *  0 * atan( 1 / (  1 + 2^24 ) )   n = 24   d_n = 1 
assign v[4'b0001] [24] = 21'h 000000;  // +0.0000000000000000 = 2^(25+1) *  0 * atan( 1 / (  1 + 2^25 ) )   n = 25   d_n = 1 
assign v[4'b0001] [25] = 21'h 000000;  // +0.0000000000000000 = 2^(26+1) *  0 * atan( 1 / (  1 + 2^26 ) )   n = 26   d_n = 1 
assign v[4'b0001] [26] = 21'h 000000;  // +0.0000000000000000 = 2^(27+1) *  0 * atan( 1 / (  1 + 2^27 ) )   n = 27   d_n = 1 
assign v[4'b0001] [27] = 21'h 000000;  // +0.0000000000000000 = 2^(28+1) *  0 * atan( 1 / (  1 + 2^28 ) )   n = 28   d_n = 1 
assign v[4'b0001] [28] = 21'h 000000;  // +0.0000000000000000 = 2^(29+1) *  0 * atan( 1 / (  1 + 2^29 ) )   n = 29   d_n = 1 
assign v[4'b0001] [29] = 21'h 000000;  // +0.0000000000000000 = 2^(30+1) *  0 * atan( 1 / (  1 + 2^30 ) )   n = 30   d_n = 1 
assign v[4'b0001] [30] = 21'h 000000;  // +0.0000000000000000 = 2^(31+1) *  0 * atan( 1 / (  1 + 2^31 ) )   n = 31   d_n = 1 
assign v[4'b0001] [31] = 21'h 000000;  // +0.0000000000000000 = 2^(32+1) *  0 * atan( 1 / (  1 + 2^32 ) )   n = 32   d_n = 1 
assign v[4'b0001] [32] = 21'h 000000;  // +0.0000000000000000 = 2^(33+1) *  0 * atan( 1 / (  1 + 2^33 ) )   n = 33   d_n = 1 
assign v[4'b0001] [33] = 21'h 000000;  // +0.0000000000000000 = 2^(34+1) *  0 * atan( 1 / (  1 + 2^34 ) )   n = 34   d_n = 1 
assign v[4'b0001] [34] = 21'h 000000;  // +0.0000000000000000 = 2^(35+1) *  0 * atan( 1 / (  1 + 2^35 ) )   n = 35   d_n = 1 
assign v[4'b0001] [35] = 21'h 000000;  // +0.0000000000000000 = 2^(36+1) *  0 * atan( 1 / (  1 + 2^36 ) )   n = 36   d_n = 1 
assign v[4'b0001] [36] = 21'h 000000;  // +0.0000000000000000 = 2^(37+1) *  0 * atan( 1 / (  1 + 2^37 ) )   n = 37   d_n = 1 
assign v[4'b0001] [37] = 21'h 000000;  // +0.0000000000000000 = 2^(38+1) *  0 * atan( 1 / (  1 + 2^38 ) )   n = 38   d_n = 1 
assign v[4'b0001] [38] = 21'h 000000;  // +0.0000000000000000 = 2^(39+1) *  0 * atan( 1 / (  1 + 2^39 ) )   n = 39   d_n = 1 
assign v[4'b0001] [39] = 21'h 000000;  // +0.0000000000000000 = 2^(40+1) *  0 * atan( 1 / (  1 + 2^40 ) )   n = 40   d_n = 1 
assign v[4'b0001] [40] = 21'h 000000;  // +0.0000000000000000 = 2^(41+1) *  0 * atan( 1 / (  1 + 2^41 ) )   n = 41   d_n = 1 
assign v[4'b0001] [41] = 21'h 000000;  // +0.0000000000000000 = 2^(42+1) *  0 * atan( 1 / (  1 + 2^42 ) )   n = 42   d_n = 1 
assign v[4'b0001] [42] = 21'h 000000;  // +0.0000000000000000 = 2^(43+1) *  0 * atan( 1 / (  1 + 2^43 ) )   n = 43   d_n = 1 
assign v[4'b0001] [43] = 21'h 000000;  // +0.0000000000000000 = 2^(44+1) *  0 * atan( 1 / (  1 + 2^44 ) )   n = 44   d_n = 1 
assign v[4'b0001] [44] = 21'h 000000;  // +0.0000000000000000 = 2^(45+1) *  0 * atan( 1 / (  1 + 2^45 ) )   n = 45   d_n = 1 
assign v[4'b0001] [45] = 21'h 000000;  // +0.0000000000000000 = 2^(46+1) *  0 * atan( 1 / (  1 + 2^46 ) )   n = 46   d_n = 1 
assign v[4'b0001] [46] = 21'h 000000;  // +0.0000000000000000 = 2^(47+1) *  0 * atan( 1 / (  1 + 2^47 ) )   n = 47   d_n = 1 
assign v[4'b0001] [47] = 21'h 000000;  // +0.0000000000000000 = 2^(48+1) *  0 * atan( 1 / (  1 + 2^48 ) )   n = 48   d_n = 1 
assign v[4'b0001] [48] = 21'h 000000;  // +0.0000000000000000 = 2^(49+1) *  0 * atan( 1 / (  1 + 2^49 ) )   n = 49   d_n = 1 
assign v[4'b0001] [49] = 21'h 000000;  // +0.0000000000000000 = 2^(50+1) *  0 * atan( 1 / (  1 + 2^50 ) )   n = 50   d_n = 1 
assign v[4'b0001] [50] = 21'h 000000;  // +0.0000000000000000 = 2^(51+1) *  0 * atan( 1 / (  1 + 2^51 ) )   n = 51   d_n = 1 
assign v[4'b0001] [51] = 21'h 000000;  // +0.0000000000000000 = 2^(52+1) *  0 * atan( 1 / (  1 + 2^52 ) )   n = 52   d_n = 1 
assign v[4'b0001] [52] = 21'h 000000;  // +0.0000000000000000 = 2^(53+1) *  0 * atan( 1 / (  1 + 2^53 ) )   n = 53   d_n = 1 
assign v[4'b0001] [53] = 21'h 000000;  // +0.0000000000000000 = 2^(54+1) *  0 * atan( 1 / (  1 + 2^54 ) )   n = 54   d_n = 1 
assign v[4'b0001] [54] = 21'h 000000;  // +0.0000000000000000 = 2^(55+1) *  0 * atan( 1 / (  1 + 2^55 ) )   n = 55   d_n = 1 
assign v[4'b0001] [55] = 21'h 000000;  // +0.0000000000000000 = 2^(56+1) *  0 * atan( 1 / (  1 + 2^56 ) )   n = 56   d_n = 1 
assign v[4'b0001] [56] = 21'h 000000;  // +0.0000000000000000 = 2^(57+1) *  0 * atan( 1 / (  1 + 2^57 ) )   n = 57   d_n = 1 
assign v[4'b0001] [57] = 21'h 000000;  // +0.0000000000000000 = 2^(58+1) *  0 * atan( 1 / (  1 + 2^58 ) )   n = 58   d_n = 1 
assign v[4'b0001] [58] = 21'h 000000;  // +0.0000000000000000 = 2^(59+1) *  0 * atan( 1 / (  1 + 2^59 ) )   n = 59   d_n = 1 
assign v[4'b0001] [59] = 21'h 000000;  // +0.0000000000000000 = 2^(60+1) *  0 * atan( 1 / (  1 + 2^60 ) )   n = 60   d_n = 1 
assign v[4'b0001] [60] = 21'h 000000;  // +0.0000000000000000 = 2^(61+1) *  0 * atan( 1 / (  1 + 2^61 ) )   n = 61   d_n = 1 
assign v[4'b0001] [61] = 21'h 000000;  // +0.0000000000000000 = 2^(62+1) *  0 * atan( 1 / (  1 + 2^62 ) )   n = 62   d_n = 1 
assign v[4'b0001] [62] = 21'h 000000;  // +0.0000000000000000 = 2^(63+1) *  0 * atan( 1 / (  1 + 2^63 ) )   n = 63   d_n = 1 
assign v[4'b0001] [63] = 21'h 000000;  // +0.0000000000000000 = 2^(64+1) *  0 * atan( 1 / (  1 + 2^64 ) )   n = 64   d_n = 1 
assign v[4'b0010] [00] = 21'h 000000;  // +0.0000000000000000 = 2^(1+1) *  0 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = -0 
assign v[4'b0010] [01] = 21'h 000000;  // +0.0000000000000000 = 2^(2+1) *  0 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = -0 
assign v[4'b0010] [02] = 21'h 000000;  // +0.0000000000000000 = 2^(3+1) *  0 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = -0 
assign v[4'b0010] [03] = 21'h 000000;  // +0.0000000000000000 = 2^(4+1) *  0 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = -0 
assign v[4'b0010] [04] = 21'h 000000;  // +0.0000000000000000 = 2^(5+1) *  0 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = -0 
assign v[4'b0010] [05] = 21'h 000000;  // +0.0000000000000000 = 2^(6+1) *  0 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = -0 
assign v[4'b0010] [06] = 21'h 000000;  // +0.0000000000000000 = 2^(7+1) *  0 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = -0 
assign v[4'b0010] [07] = 21'h 000000;  // +0.0000000000000000 = 2^(8+1) *  0 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = -0 
assign v[4'b0010] [08] = 21'h 000000;  // +0.0000000000000000 = 2^(9+1) *  0 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = -0 
assign v[4'b0010] [09] = 21'h 000000;  // +0.0000000000000000 = 2^(10+1) *  0 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = -0 
assign v[4'b0010] [10] = 21'h 000000;  // +0.0000000000000000 = 2^(11+1) *  0 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = -0 
assign v[4'b0010] [11] = 21'h 000000;  // +0.0000000000000000 = 2^(12+1) *  0 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = -0 
assign v[4'b0010] [12] = 21'h 000000;  // +0.0000000000000000 = 2^(13+1) *  0 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = -0 
assign v[4'b0010] [13] = 21'h 000000;  // +0.0000000000000000 = 2^(14+1) *  0 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = -0 
assign v[4'b0010] [14] = 21'h 000000;  // +0.0000000000000000 = 2^(15+1) *  0 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = -0 
assign v[4'b0010] [15] = 21'h 000000;  // +0.0000000000000000 = 2^(16+1) *  0 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = -0 
assign v[4'b0010] [16] = 21'h 000000;  // +0.0000000000000000 = 2^(17+1) *  0 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = -0 
assign v[4'b0010] [17] = 21'h 000000;  // +0.0000000000000000 = 2^(18+1) *  0 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = -0 
assign v[4'b0010] [18] = 21'h 000000;  // +0.0000000000000000 = 2^(19+1) *  0 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = -0 
assign v[4'b0010] [19] = 21'h 000000;  // +0.0000000000000000 = 2^(20+1) *  0 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = -0 
assign v[4'b0010] [20] = 21'h 000000;  // +0.0000000000000000 = 2^(21+1) *  0 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = -0 
assign v[4'b0010] [21] = 21'h 000000;  // +0.0000000000000000 = 2^(22+1) *  0 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = -0 
assign v[4'b0010] [22] = 21'h 000000;  // +0.0000000000000000 = 2^(23+1) *  0 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = -0 
assign v[4'b0010] [23] = 21'h 000000;  // +0.0000000000000000 = 2^(24+1) *  0 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = -0 
assign v[4'b0010] [24] = 21'h 000000;  // +0.0000000000000000 = 2^(25+1) *  0 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = -0 
assign v[4'b0010] [25] = 21'h 000000;  // +0.0000000000000000 = 2^(26+1) *  0 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = -0 
assign v[4'b0010] [26] = 21'h 000000;  // +0.0000000000000000 = 2^(27+1) *  0 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = -0 
assign v[4'b0010] [27] = 21'h 000000;  // +0.0000000000000000 = 2^(28+1) *  0 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = -0 
assign v[4'b0010] [28] = 21'h 000000;  // +0.0000000000000000 = 2^(29+1) *  0 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = -0 
assign v[4'b0010] [29] = 21'h 000000;  // +0.0000000000000000 = 2^(30+1) *  0 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = -0 
assign v[4'b0010] [30] = 21'h 000000;  // +0.0000000000000000 = 2^(31+1) *  0 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = -0 
assign v[4'b0010] [31] = 21'h 000000;  // +0.0000000000000000 = 2^(32+1) *  0 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = -0 
assign v[4'b0010] [32] = 21'h 000000;  // +0.0000000000000000 = 2^(33+1) *  0 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = -0 
assign v[4'b0010] [33] = 21'h 000000;  // +0.0000000000000000 = 2^(34+1) *  0 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = -0 
assign v[4'b0010] [34] = 21'h 000000;  // +0.0000000000000000 = 2^(35+1) *  0 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = -0 
assign v[4'b0010] [35] = 21'h 000000;  // +0.0000000000000000 = 2^(36+1) *  0 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = -0 
assign v[4'b0010] [36] = 21'h 000000;  // +0.0000000000000000 = 2^(37+1) *  0 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = -0 
assign v[4'b0010] [37] = 21'h 000000;  // +0.0000000000000000 = 2^(38+1) *  0 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = -0 
assign v[4'b0010] [38] = 21'h 000000;  // +0.0000000000000000 = 2^(39+1) *  0 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = -0 
assign v[4'b0010] [39] = 21'h 000000;  // +0.0000000000000000 = 2^(40+1) *  0 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = -0 
assign v[4'b0010] [40] = 21'h 000000;  // +0.0000000000000000 = 2^(41+1) *  0 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = -0 
assign v[4'b0010] [41] = 21'h 000000;  // +0.0000000000000000 = 2^(42+1) *  0 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = -0 
assign v[4'b0010] [42] = 21'h 000000;  // +0.0000000000000000 = 2^(43+1) *  0 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = -0 
assign v[4'b0010] [43] = 21'h 000000;  // +0.0000000000000000 = 2^(44+1) *  0 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = -0 
assign v[4'b0010] [44] = 21'h 000000;  // +0.0000000000000000 = 2^(45+1) *  0 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = -0 
assign v[4'b0010] [45] = 21'h 000000;  // +0.0000000000000000 = 2^(46+1) *  0 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = -0 
assign v[4'b0010] [46] = 21'h 000000;  // +0.0000000000000000 = 2^(47+1) *  0 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = -0 
assign v[4'b0010] [47] = 21'h 000000;  // +0.0000000000000000 = 2^(48+1) *  0 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = -0 
assign v[4'b0010] [48] = 21'h 000000;  // +0.0000000000000000 = 2^(49+1) *  0 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = -0 
assign v[4'b0010] [49] = 21'h 000000;  // +0.0000000000000000 = 2^(50+1) *  0 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = -0 
assign v[4'b0010] [50] = 21'h 000000;  // +0.0000000000000000 = 2^(51+1) *  0 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = -0 
assign v[4'b0010] [51] = 21'h 000000;  // +0.0000000000000000 = 2^(52+1) *  0 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = -0 
assign v[4'b0010] [52] = 21'h 000000;  // +0.0000000000000000 = 2^(53+1) *  0 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = -0 
assign v[4'b0010] [53] = 21'h 000000;  // +0.0000000000000000 = 2^(54+1) *  0 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = -0 
assign v[4'b0010] [54] = 21'h 000000;  // +0.0000000000000000 = 2^(55+1) *  0 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = -0 
assign v[4'b0010] [55] = 21'h 000000;  // +0.0000000000000000 = 2^(56+1) *  0 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = -0 
assign v[4'b0010] [56] = 21'h 000000;  // +0.0000000000000000 = 2^(57+1) *  0 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = -0 
assign v[4'b0010] [57] = 21'h 000000;  // +0.0000000000000000 = 2^(58+1) *  0 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = -0 
assign v[4'b0010] [58] = 21'h 000000;  // +0.0000000000000000 = 2^(59+1) *  0 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = -0 
assign v[4'b0010] [59] = 21'h 000000;  // +0.0000000000000000 = 2^(60+1) *  0 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = -0 
assign v[4'b0010] [60] = 21'h 000000;  // +0.0000000000000000 = 2^(61+1) *  0 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = -0 
assign v[4'b0010] [61] = 21'h 000000;  // +0.0000000000000000 = 2^(62+1) *  0 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = -0 
assign v[4'b0010] [62] = 21'h 000000;  // +0.0000000000000000 = 2^(63+1) *  0 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = -0 
assign v[4'b0010] [63] = 21'h 000000;  // +0.0000000000000000 = 2^(64+1) *  0 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = -0 
assign v[4'b0011] [00] = 21'h 000000;  // -0.0000000000000000 = 2^(1+1) *  0 * atan( 1 / ( -1 + 2^1 ) )   n =  1   d_n = -1 
assign v[4'b0011] [01] = 21'h 000000;  // -0.0000000000000000 = 2^(2+1) *  0 * atan( 1 / ( -1 + 2^2 ) )   n =  2   d_n = -1 
assign v[4'b0011] [02] = 21'h 000000;  // -0.0000000000000000 = 2^(3+1) *  0 * atan( 1 / ( -1 + 2^3 ) )   n =  3   d_n = -1 
assign v[4'b0011] [03] = 21'h 000000;  // -0.0000000000000000 = 2^(4+1) *  0 * atan( 1 / ( -1 + 2^4 ) )   n =  4   d_n = -1 
assign v[4'b0011] [04] = 21'h 000000;  // -0.0000000000000000 = 2^(5+1) *  0 * atan( 1 / ( -1 + 2^5 ) )   n =  5   d_n = -1 
assign v[4'b0011] [05] = 21'h 000000;  // -0.0000000000000000 = 2^(6+1) *  0 * atan( 1 / ( -1 + 2^6 ) )   n =  6   d_n = -1 
assign v[4'b0011] [06] = 21'h 000000;  // -0.0000000000000000 = 2^(7+1) *  0 * atan( 1 / ( -1 + 2^7 ) )   n =  7   d_n = -1 
assign v[4'b0011] [07] = 21'h 000000;  // -0.0000000000000000 = 2^(8+1) *  0 * atan( 1 / ( -1 + 2^8 ) )   n =  8   d_n = -1 
assign v[4'b0011] [08] = 21'h 000000;  // -0.0000000000000000 = 2^(9+1) *  0 * atan( 1 / ( -1 + 2^9 ) )   n =  9   d_n = -1 
assign v[4'b0011] [09] = 21'h 000000;  // -0.0000000000000000 = 2^(10+1) *  0 * atan( 1 / ( -1 + 2^10 ) )   n = 10   d_n = -1 
assign v[4'b0011] [10] = 21'h 000000;  // -0.0000000000000000 = 2^(11+1) *  0 * atan( 1 / ( -1 + 2^11 ) )   n = 11   d_n = -1 
assign v[4'b0011] [11] = 21'h 000000;  // -0.0000000000000000 = 2^(12+1) *  0 * atan( 1 / ( -1 + 2^12 ) )   n = 12   d_n = -1 
assign v[4'b0011] [12] = 21'h 000000;  // -0.0000000000000000 = 2^(13+1) *  0 * atan( 1 / ( -1 + 2^13 ) )   n = 13   d_n = -1 
assign v[4'b0011] [13] = 21'h 000000;  // -0.0000000000000000 = 2^(14+1) *  0 * atan( 1 / ( -1 + 2^14 ) )   n = 14   d_n = -1 
assign v[4'b0011] [14] = 21'h 000000;  // -0.0000000000000000 = 2^(15+1) *  0 * atan( 1 / ( -1 + 2^15 ) )   n = 15   d_n = -1 
assign v[4'b0011] [15] = 21'h 000000;  // -0.0000000000000000 = 2^(16+1) *  0 * atan( 1 / ( -1 + 2^16 ) )   n = 16   d_n = -1 
assign v[4'b0011] [16] = 21'h 000000;  // -0.0000000000000000 = 2^(17+1) *  0 * atan( 1 / ( -1 + 2^17 ) )   n = 17   d_n = -1 
assign v[4'b0011] [17] = 21'h 000000;  // -0.0000000000000000 = 2^(18+1) *  0 * atan( 1 / ( -1 + 2^18 ) )   n = 18   d_n = -1 
assign v[4'b0011] [18] = 21'h 000000;  // -0.0000000000000000 = 2^(19+1) *  0 * atan( 1 / ( -1 + 2^19 ) )   n = 19   d_n = -1 
assign v[4'b0011] [19] = 21'h 000000;  // -0.0000000000000000 = 2^(20+1) *  0 * atan( 1 / ( -1 + 2^20 ) )   n = 20   d_n = -1 
assign v[4'b0011] [20] = 21'h 000000;  // -0.0000000000000000 = 2^(21+1) *  0 * atan( 1 / ( -1 + 2^21 ) )   n = 21   d_n = -1 
assign v[4'b0011] [21] = 21'h 000000;  // -0.0000000000000000 = 2^(22+1) *  0 * atan( 1 / ( -1 + 2^22 ) )   n = 22   d_n = -1 
assign v[4'b0011] [22] = 21'h 000000;  // -0.0000000000000000 = 2^(23+1) *  0 * atan( 1 / ( -1 + 2^23 ) )   n = 23   d_n = -1 
assign v[4'b0011] [23] = 21'h 000000;  // -0.0000000000000000 = 2^(24+1) *  0 * atan( 1 / ( -1 + 2^24 ) )   n = 24   d_n = -1 
assign v[4'b0011] [24] = 21'h 000000;  // -0.0000000000000000 = 2^(25+1) *  0 * atan( 1 / ( -1 + 2^25 ) )   n = 25   d_n = -1 
assign v[4'b0011] [25] = 21'h 000000;  // -0.0000000000000000 = 2^(26+1) *  0 * atan( 1 / ( -1 + 2^26 ) )   n = 26   d_n = -1 
assign v[4'b0011] [26] = 21'h 000000;  // -0.0000000000000000 = 2^(27+1) *  0 * atan( 1 / ( -1 + 2^27 ) )   n = 27   d_n = -1 
assign v[4'b0011] [27] = 21'h 000000;  // -0.0000000000000000 = 2^(28+1) *  0 * atan( 1 / ( -1 + 2^28 ) )   n = 28   d_n = -1 
assign v[4'b0011] [28] = 21'h 000000;  // -0.0000000000000000 = 2^(29+1) *  0 * atan( 1 / ( -1 + 2^29 ) )   n = 29   d_n = -1 
assign v[4'b0011] [29] = 21'h 000000;  // -0.0000000000000000 = 2^(30+1) *  0 * atan( 1 / ( -1 + 2^30 ) )   n = 30   d_n = -1 
assign v[4'b0011] [30] = 21'h 000000;  // -0.0000000000000000 = 2^(31+1) *  0 * atan( 1 / ( -1 + 2^31 ) )   n = 31   d_n = -1 
assign v[4'b0011] [31] = 21'h 000000;  // -0.0000000000000000 = 2^(32+1) *  0 * atan( 1 / ( -1 + 2^32 ) )   n = 32   d_n = -1 
assign v[4'b0011] [32] = 21'h 000000;  // -0.0000000000000000 = 2^(33+1) *  0 * atan( 1 / ( -1 + 2^33 ) )   n = 33   d_n = -1 
assign v[4'b0011] [33] = 21'h 000000;  // -0.0000000000000000 = 2^(34+1) *  0 * atan( 1 / ( -1 + 2^34 ) )   n = 34   d_n = -1 
assign v[4'b0011] [34] = 21'h 000000;  // -0.0000000000000000 = 2^(35+1) *  0 * atan( 1 / ( -1 + 2^35 ) )   n = 35   d_n = -1 
assign v[4'b0011] [35] = 21'h 000000;  // -0.0000000000000000 = 2^(36+1) *  0 * atan( 1 / ( -1 + 2^36 ) )   n = 36   d_n = -1 
assign v[4'b0011] [36] = 21'h 000000;  // -0.0000000000000000 = 2^(37+1) *  0 * atan( 1 / ( -1 + 2^37 ) )   n = 37   d_n = -1 
assign v[4'b0011] [37] = 21'h 000000;  // -0.0000000000000000 = 2^(38+1) *  0 * atan( 1 / ( -1 + 2^38 ) )   n = 38   d_n = -1 
assign v[4'b0011] [38] = 21'h 000000;  // -0.0000000000000000 = 2^(39+1) *  0 * atan( 1 / ( -1 + 2^39 ) )   n = 39   d_n = -1 
assign v[4'b0011] [39] = 21'h 000000;  // -0.0000000000000000 = 2^(40+1) *  0 * atan( 1 / ( -1 + 2^40 ) )   n = 40   d_n = -1 
assign v[4'b0011] [40] = 21'h 000000;  // -0.0000000000000000 = 2^(41+1) *  0 * atan( 1 / ( -1 + 2^41 ) )   n = 41   d_n = -1 
assign v[4'b0011] [41] = 21'h 000000;  // -0.0000000000000000 = 2^(42+1) *  0 * atan( 1 / ( -1 + 2^42 ) )   n = 42   d_n = -1 
assign v[4'b0011] [42] = 21'h 000000;  // -0.0000000000000000 = 2^(43+1) *  0 * atan( 1 / ( -1 + 2^43 ) )   n = 43   d_n = -1 
assign v[4'b0011] [43] = 21'h 000000;  // -0.0000000000000000 = 2^(44+1) *  0 * atan( 1 / ( -1 + 2^44 ) )   n = 44   d_n = -1 
assign v[4'b0011] [44] = 21'h 000000;  // -0.0000000000000000 = 2^(45+1) *  0 * atan( 1 / ( -1 + 2^45 ) )   n = 45   d_n = -1 
assign v[4'b0011] [45] = 21'h 000000;  // -0.0000000000000000 = 2^(46+1) *  0 * atan( 1 / ( -1 + 2^46 ) )   n = 46   d_n = -1 
assign v[4'b0011] [46] = 21'h 000000;  // -0.0000000000000000 = 2^(47+1) *  0 * atan( 1 / ( -1 + 2^47 ) )   n = 47   d_n = -1 
assign v[4'b0011] [47] = 21'h 000000;  // -0.0000000000000000 = 2^(48+1) *  0 * atan( 1 / ( -1 + 2^48 ) )   n = 48   d_n = -1 
assign v[4'b0011] [48] = 21'h 000000;  // -0.0000000000000000 = 2^(49+1) *  0 * atan( 1 / ( -1 + 2^49 ) )   n = 49   d_n = -1 
assign v[4'b0011] [49] = 21'h 000000;  // -0.0000000000000000 = 2^(50+1) *  0 * atan( 1 / ( -1 + 2^50 ) )   n = 50   d_n = -1 
assign v[4'b0011] [50] = 21'h 000000;  // -0.0000000000000000 = 2^(51+1) *  0 * atan( 1 / ( -1 + 2^51 ) )   n = 51   d_n = -1 
assign v[4'b0011] [51] = 21'h 000000;  // -0.0000000000000000 = 2^(52+1) *  0 * atan( 1 / ( -1 + 2^52 ) )   n = 52   d_n = -1 
assign v[4'b0011] [52] = 21'h 000000;  // -0.0000000000000000 = 2^(53+1) *  0 * atan( 1 / ( -1 + 2^53 ) )   n = 53   d_n = -1 
assign v[4'b0011] [53] = 21'h 000000;  // -0.0000000000000000 = 2^(54+1) *  0 * atan( 1 / ( -1 + 2^54 ) )   n = 54   d_n = -1 
assign v[4'b0011] [54] = 21'h 000000;  // -0.0000000000000000 = 2^(55+1) *  0 * atan( 1 / ( -1 + 2^55 ) )   n = 55   d_n = -1 
assign v[4'b0011] [55] = 21'h 000000;  // -0.0000000000000000 = 2^(56+1) *  0 * atan( 1 / ( -1 + 2^56 ) )   n = 56   d_n = -1 
assign v[4'b0011] [56] = 21'h 000000;  // -0.0000000000000000 = 2^(57+1) *  0 * atan( 1 / ( -1 + 2^57 ) )   n = 57   d_n = -1 
assign v[4'b0011] [57] = 21'h 000000;  // -0.0000000000000000 = 2^(58+1) *  0 * atan( 1 / ( -1 + 2^58 ) )   n = 58   d_n = -1 
assign v[4'b0011] [58] = 21'h 000000;  // -0.0000000000000000 = 2^(59+1) *  0 * atan( 1 / ( -1 + 2^59 ) )   n = 59   d_n = -1 
assign v[4'b0011] [59] = 21'h 000000;  // -0.0000000000000000 = 2^(60+1) *  0 * atan( 1 / ( -1 + 2^60 ) )   n = 60   d_n = -1 
assign v[4'b0011] [60] = 21'h 000000;  // -0.0000000000000000 = 2^(61+1) *  0 * atan( 1 / ( -1 + 2^61 ) )   n = 61   d_n = -1 
assign v[4'b0011] [61] = 21'h 000000;  // -0.0000000000000000 = 2^(62+1) *  0 * atan( 1 / ( -1 + 2^62 ) )   n = 62   d_n = -1 
assign v[4'b0011] [62] = 21'h 000000;  // -0.0000000000000000 = 2^(63+1) *  0 * atan( 1 / ( -1 + 2^63 ) )   n = 63   d_n = -1 
assign v[4'b0011] [63] = 21'h 000000;  // -0.0000000000000000 = 2^(64+1) *  0 * atan( 1 / ( -1 + 2^64 ) )   n = 64   d_n = -1 
assign v[4'b0100] [00] = 21'h 00076B;  // +1.8545904360032244 = 2^(1+1) *  1 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = 0+1i 
assign v[4'b0100] [01] = 21'h 0007D6;  // +1.9598293050149131 = 2^(2+1) *  1 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = 0+1i 
assign v[4'b0100] [02] = 21'h 0007F5;  // +1.9896799127481830 = 2^(3+1) *  1 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = 0+1i 
assign v[4'b0100] [03] = 21'h 0007FD;  // +1.9974019198706352 = 2^(4+1) *  1 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = 0+1i 
assign v[4'b0100] [04] = 21'h 0007FF;  // +1.9993493395371698 = 2^(5+1) *  1 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = 0+1i 
assign v[4'b0100] [05] = 21'h 0007FF;  // +1.9998372634210344 = 2^(6+1) *  1 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = 0+1i 
assign v[4'b0100] [06] = 21'h 0007FF;  // +1.9999593113858845 = 2^(7+1) *  1 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = 0+1i 
assign v[4'b0100] [07] = 21'h 0007FF;  // +1.9999898275670895 = 2^(8+1) *  1 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = 0+1i 
assign v[4'b0100] [08] = 21'h 0007FF;  // +1.9999974568743104 = 2^(9+1) *  1 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = 0+1i 
assign v[4'b0100] [09] = 21'h 0007FF;  // +1.9999993642174863 = 2^(10+1) *  1 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = 0+1i 
assign v[4'b0100] [10] = 21'h 0007FF;  // +1.9999998410543034 = 2^(11+1) *  1 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = 0+1i 
assign v[4'b0100] [11] = 21'h 0007FF;  // +1.9999999602635716 = 2^(12+1) *  1 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = 0+1i 
assign v[4'b0100] [12] = 21'h 0007FF;  // +1.9999999900658927 = 2^(13+1) *  1 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = 0+1i 
assign v[4'b0100] [13] = 21'h 0007FF;  // +1.9999999975164731 = 2^(14+1) *  1 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = 0+1i 
assign v[4'b0100] [14] = 21'h 0007FF;  // +1.9999999993791182 = 2^(15+1) *  1 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = 0+1i 
assign v[4'b0100] [15] = 21'h 0007FF;  // +1.9999999998447795 = 2^(16+1) *  1 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = 0+1i 
assign v[4'b0100] [16] = 21'h 0007FF;  // +1.9999999999611948 = 2^(17+1) *  1 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = 0+1i 
assign v[4'b0100] [17] = 21'h 0007FF;  // +1.9999999999902986 = 2^(18+1) *  1 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = 0+1i 
assign v[4'b0100] [18] = 21'h 0007FF;  // +1.9999999999975746 = 2^(19+1) *  1 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = 0+1i 
assign v[4'b0100] [19] = 21'h 0007FF;  // +1.9999999999993936 = 2^(20+1) *  1 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = 0+1i 
assign v[4'b0100] [20] = 21'h 0007FF;  // +1.9999999999998483 = 2^(21+1) *  1 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = 0+1i 
assign v[4'b0100] [21] = 21'h 0007FF;  // +1.9999999999999620 = 2^(22+1) *  1 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = 0+1i 
assign v[4'b0100] [22] = 21'h 0007FF;  // +1.9999999999999905 = 2^(23+1) *  1 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = 0+1i 
assign v[4'b0100] [23] = 21'h 0007FF;  // +1.9999999999999976 = 2^(24+1) *  1 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = 0+1i 
assign v[4'b0100] [24] = 21'h 0007FF;  // +1.9999999999999993 = 2^(25+1) *  1 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = 0+1i 
assign v[4'b0100] [25] = 21'h 0007FF;  // +1.9999999999999998 = 2^(26+1) *  1 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = 0+1i 
assign v[4'b0100] [26] = 21'h 000800;  // +2.0000000000000000 = 2^(27+1) *  1 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = 0+1i 
assign v[4'b0100] [27] = 21'h 000800;  // +2.0000000000000000 = 2^(28+1) *  1 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = 0+1i 
assign v[4'b0100] [28] = 21'h 000800;  // +2.0000000000000000 = 2^(29+1) *  1 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = 0+1i 
assign v[4'b0100] [29] = 21'h 000800;  // +2.0000000000000000 = 2^(30+1) *  1 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = 0+1i 
assign v[4'b0100] [30] = 21'h 000800;  // +2.0000000000000000 = 2^(31+1) *  1 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = 0+1i 
assign v[4'b0100] [31] = 21'h 000800;  // +2.0000000000000000 = 2^(32+1) *  1 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = 0+1i 
assign v[4'b0100] [32] = 21'h 000800;  // +2.0000000000000000 = 2^(33+1) *  1 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = 0+1i 
assign v[4'b0100] [33] = 21'h 000800;  // +2.0000000000000000 = 2^(34+1) *  1 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = 0+1i 
assign v[4'b0100] [34] = 21'h 000800;  // +2.0000000000000000 = 2^(35+1) *  1 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = 0+1i 
assign v[4'b0100] [35] = 21'h 000800;  // +2.0000000000000000 = 2^(36+1) *  1 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = 0+1i 
assign v[4'b0100] [36] = 21'h 000800;  // +2.0000000000000000 = 2^(37+1) *  1 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = 0+1i 
assign v[4'b0100] [37] = 21'h 000800;  // +2.0000000000000000 = 2^(38+1) *  1 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = 0+1i 
assign v[4'b0100] [38] = 21'h 000800;  // +2.0000000000000000 = 2^(39+1) *  1 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = 0+1i 
assign v[4'b0100] [39] = 21'h 000800;  // +2.0000000000000000 = 2^(40+1) *  1 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = 0+1i 
assign v[4'b0100] [40] = 21'h 000800;  // +2.0000000000000000 = 2^(41+1) *  1 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = 0+1i 
assign v[4'b0100] [41] = 21'h 000800;  // +2.0000000000000000 = 2^(42+1) *  1 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = 0+1i 
assign v[4'b0100] [42] = 21'h 000800;  // +2.0000000000000000 = 2^(43+1) *  1 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = 0+1i 
assign v[4'b0100] [43] = 21'h 000800;  // +2.0000000000000000 = 2^(44+1) *  1 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = 0+1i 
assign v[4'b0100] [44] = 21'h 000800;  // +2.0000000000000000 = 2^(45+1) *  1 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = 0+1i 
assign v[4'b0100] [45] = 21'h 000800;  // +2.0000000000000000 = 2^(46+1) *  1 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = 0+1i 
assign v[4'b0100] [46] = 21'h 000800;  // +2.0000000000000000 = 2^(47+1) *  1 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = 0+1i 
assign v[4'b0100] [47] = 21'h 000800;  // +2.0000000000000000 = 2^(48+1) *  1 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = 0+1i 
assign v[4'b0100] [48] = 21'h 000800;  // +2.0000000000000000 = 2^(49+1) *  1 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = 0+1i 
assign v[4'b0100] [49] = 21'h 000800;  // +2.0000000000000000 = 2^(50+1) *  1 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = 0+1i 
assign v[4'b0100] [50] = 21'h 000800;  // +2.0000000000000000 = 2^(51+1) *  1 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = 0+1i 
assign v[4'b0100] [51] = 21'h 000800;  // +2.0000000000000000 = 2^(52+1) *  1 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = 0+1i 
assign v[4'b0100] [52] = 21'h 000800;  // +2.0000000000000000 = 2^(53+1) *  1 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = 0+1i 
assign v[4'b0100] [53] = 21'h 000800;  // +2.0000000000000000 = 2^(54+1) *  1 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = 0+1i 
assign v[4'b0100] [54] = 21'h 000800;  // +2.0000000000000000 = 2^(55+1) *  1 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = 0+1i 
assign v[4'b0100] [55] = 21'h 000800;  // +2.0000000000000000 = 2^(56+1) *  1 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = 0+1i 
assign v[4'b0100] [56] = 21'h 000800;  // +2.0000000000000000 = 2^(57+1) *  1 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = 0+1i 
assign v[4'b0100] [57] = 21'h 000800;  // +2.0000000000000000 = 2^(58+1) *  1 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = 0+1i 
assign v[4'b0100] [58] = 21'h 000800;  // +2.0000000000000000 = 2^(59+1) *  1 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = 0+1i 
assign v[4'b0100] [59] = 21'h 000800;  // +2.0000000000000000 = 2^(60+1) *  1 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = 0+1i 
assign v[4'b0100] [60] = 21'h 000800;  // +2.0000000000000000 = 2^(61+1) *  1 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = 0+1i 
assign v[4'b0100] [61] = 21'h 000800;  // +2.0000000000000000 = 2^(62+1) *  1 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = 0+1i 
assign v[4'b0100] [62] = 21'h 000800;  // +2.0000000000000000 = 2^(63+1) *  1 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = 0+1i 
assign v[4'b0100] [63] = 21'h 000800;  // +2.0000000000000000 = 2^(64+1) *  1 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = 0+1i 
assign v[4'b0101] [00] = 21'h 000525;  // +1.2870022175865687 = 2^(1+1) *  1 * atan( 1 / (  1 + 2^1 ) )   n =  1   d_n = 1+1i 
assign v[4'b0101] [01] = 21'h 000651;  // +1.5791644787990460 = 2^(2+1) *  1 * atan( 1 / (  1 + 2^2 ) )   n =  2   d_n = 1+1i 
assign v[4'b0101] [02] = 21'h 000715;  // +1.7705155387823304 = 2^(3+1) *  1 * atan( 1 / (  1 + 2^3 ) )   n =  3   d_n = 1+1i 
assign v[4'b0101] [03] = 21'h 000785;  // +1.8801863269031263 = 2^(4+1) *  1 * atan( 1 / (  1 + 2^4 ) )   n =  4   d_n = 1+1i 
assign v[4'b0101] [04] = 21'h 0007C1;  // +1.9388006348016065 = 2^(5+1) *  1 * atan( 1 / (  1 + 2^5 ) )   n =  5   d_n = 1+1i 
assign v[4'b0101] [05] = 21'h 0007E0;  // +1.9690754279161793 = 2^(6+1) *  1 * atan( 1 / (  1 + 2^6 ) )   n =  6   d_n = 1+1i 
assign v[4'b0101] [06] = 21'h 0007F0;  // +1.9844563743249595 = 2^(7+1) *  1 * atan( 1 / (  1 + 2^7 ) )   n =  7   d_n = 1+1i 
assign v[4'b0101] [07] = 21'h 0007F8;  // +1.9922078446819715 = 2^(8+1) *  1 * atan( 1 / (  1 + 2^8 ) )   n =  8   d_n = 1+1i 
assign v[4'b0101] [08] = 21'h 0007FC;  // +1.9960988362398133 = 2^(9+1) *  1 * atan( 1 / (  1 + 2^9 ) )   n =  9   d_n = 1+1i 
assign v[4'b0101] [09] = 21'h 0007FE;  // +1.9980481465643023 = 2^(10+1) *  1 * atan( 1 / (  1 + 2^10 ) )   n = 10   d_n = 1+1i 
assign v[4'b0101] [10] = 21'h 0007FF;  // +1.9990237553913479 = 2^(11+1) *  1 * atan( 1 / (  1 + 2^11 ) )   n = 11   d_n = 1+1i 
assign v[4'b0101] [11] = 21'h 0007FF;  // +1.9995117982228541 = 2^(12+1) *  1 * atan( 1 / (  1 + 2^12 ) )   n = 12   d_n = 1+1i 
assign v[4'b0101] [12] = 21'h 0007FF;  // +1.9997558792432146 = 2^(13+1) *  1 * atan( 1 / (  1 + 2^13 ) )   n = 13   d_n = 1+1i 
assign v[4'b0101] [13] = 21'h 0007FF;  // +1.9998779346545537 = 2^(14+1) *  1 * atan( 1 / (  1 + 2^14 ) )   n = 14   d_n = 1+1i 
assign v[4'b0101] [14] = 21'h 0007FF;  // +1.9999389660855134 = 2^(15+1) *  1 * atan( 1 / (  1 + 2^15 ) )   n = 15   d_n = 1+1i 
assign v[4'b0101] [15] = 21'h 0007FF;  // +1.9999694827323158 = 2^(16+1) *  1 * atan( 1 / (  1 + 2^16 ) )   n = 16   d_n = 1+1i 
assign v[4'b0101] [16] = 21'h 0007FF;  // +1.9999847412885476 = 2^(17+1) *  1 * atan( 1 / (  1 + 2^17 ) )   n = 17   d_n = 1+1i 
assign v[4'b0101] [17] = 21'h 0007FF;  // +1.9999923706248712 = 2^(18+1) *  1 * atan( 1 / (  1 + 2^18 ) )   n = 18   d_n = 1+1i 
assign v[4'b0101] [18] = 21'h 0007FF;  // +1.9999961853075849 = 2^(19+1) *  1 * atan( 1 / (  1 + 2^19 ) )   n = 19   d_n = 1+1i 
assign v[4'b0101] [19] = 21'h 0007FF;  // +1.9999980926525798 = 2^(20+1) *  1 * atan( 1 / (  1 + 2^20 ) )   n = 20   d_n = 1+1i 
assign v[4'b0101] [20] = 21'h 0007FF;  // +1.9999990463259867 = 2^(21+1) *  1 * atan( 1 / (  1 + 2^21 ) )   n = 21   d_n = 1+1i 
assign v[4'b0101] [21] = 21'h 0007FF;  // +1.9999995231629175 = 2^(22+1) *  1 * atan( 1 / (  1 + 2^22 ) )   n = 22   d_n = 1+1i 
assign v[4'b0101] [22] = 21'h 0007FF;  // +1.9999997615814398 = 2^(23+1) *  1 * atan( 1 / (  1 + 2^23 ) )   n = 23   d_n = 1+1i 
assign v[4'b0101] [23] = 21'h 0007FF;  // +1.9999998807907151 = 2^(24+1) *  1 * atan( 1 / (  1 + 2^24 ) )   n = 24   d_n = 1+1i 
assign v[4'b0101] [24] = 21'h 0007FF;  // +1.9999999403953563 = 2^(25+1) *  1 * atan( 1 / (  1 + 2^25 ) )   n = 25   d_n = 1+1i 
assign v[4'b0101] [25] = 21'h 0007FF;  // +1.9999999701976778 = 2^(26+1) *  1 * atan( 1 / (  1 + 2^26 ) )   n = 26   d_n = 1+1i 
assign v[4'b0101] [26] = 21'h 0007FF;  // +1.9999999850988388 = 2^(27+1) *  1 * atan( 1 / (  1 + 2^27 ) )   n = 27   d_n = 1+1i 
assign v[4'b0101] [27] = 21'h 0007FF;  // +1.9999999925494194 = 2^(28+1) *  1 * atan( 1 / (  1 + 2^28 ) )   n = 28   d_n = 1+1i 
assign v[4'b0101] [28] = 21'h 0007FF;  // +1.9999999962747097 = 2^(29+1) *  1 * atan( 1 / (  1 + 2^29 ) )   n = 29   d_n = 1+1i 
assign v[4'b0101] [29] = 21'h 0007FF;  // +1.9999999981373549 = 2^(30+1) *  1 * atan( 1 / (  1 + 2^30 ) )   n = 30   d_n = 1+1i 
assign v[4'b0101] [30] = 21'h 0007FF;  // +1.9999999990686774 = 2^(31+1) *  1 * atan( 1 / (  1 + 2^31 ) )   n = 31   d_n = 1+1i 
assign v[4'b0101] [31] = 21'h 0007FF;  // +1.9999999995343387 = 2^(32+1) *  1 * atan( 1 / (  1 + 2^32 ) )   n = 32   d_n = 1+1i 
assign v[4'b0101] [32] = 21'h 0007FF;  // +1.9999999997671694 = 2^(33+1) *  1 * atan( 1 / (  1 + 2^33 ) )   n = 33   d_n = 1+1i 
assign v[4'b0101] [33] = 21'h 0007FF;  // +1.9999999998835847 = 2^(34+1) *  1 * atan( 1 / (  1 + 2^34 ) )   n = 34   d_n = 1+1i 
assign v[4'b0101] [34] = 21'h 0007FF;  // +1.9999999999417923 = 2^(35+1) *  1 * atan( 1 / (  1 + 2^35 ) )   n = 35   d_n = 1+1i 
assign v[4'b0101] [35] = 21'h 0007FF;  // +1.9999999999708962 = 2^(36+1) *  1 * atan( 1 / (  1 + 2^36 ) )   n = 36   d_n = 1+1i 
assign v[4'b0101] [36] = 21'h 0007FF;  // +1.9999999999854481 = 2^(37+1) *  1 * atan( 1 / (  1 + 2^37 ) )   n = 37   d_n = 1+1i 
assign v[4'b0101] [37] = 21'h 0007FF;  // +1.9999999999927240 = 2^(38+1) *  1 * atan( 1 / (  1 + 2^38 ) )   n = 38   d_n = 1+1i 
assign v[4'b0101] [38] = 21'h 0007FF;  // +1.9999999999963620 = 2^(39+1) *  1 * atan( 1 / (  1 + 2^39 ) )   n = 39   d_n = 1+1i 
assign v[4'b0101] [39] = 21'h 0007FF;  // +1.9999999999981810 = 2^(40+1) *  1 * atan( 1 / (  1 + 2^40 ) )   n = 40   d_n = 1+1i 
assign v[4'b0101] [40] = 21'h 0007FF;  // +1.9999999999990905 = 2^(41+1) *  1 * atan( 1 / (  1 + 2^41 ) )   n = 41   d_n = 1+1i 
assign v[4'b0101] [41] = 21'h 0007FF;  // +1.9999999999995453 = 2^(42+1) *  1 * atan( 1 / (  1 + 2^42 ) )   n = 42   d_n = 1+1i 
assign v[4'b0101] [42] = 21'h 0007FF;  // +1.9999999999997726 = 2^(43+1) *  1 * atan( 1 / (  1 + 2^43 ) )   n = 43   d_n = 1+1i 
assign v[4'b0101] [43] = 21'h 0007FF;  // +1.9999999999998863 = 2^(44+1) *  1 * atan( 1 / (  1 + 2^44 ) )   n = 44   d_n = 1+1i 
assign v[4'b0101] [44] = 21'h 0007FF;  // +1.9999999999999432 = 2^(45+1) *  1 * atan( 1 / (  1 + 2^45 ) )   n = 45   d_n = 1+1i 
assign v[4'b0101] [45] = 21'h 0007FF;  // +1.9999999999999716 = 2^(46+1) *  1 * atan( 1 / (  1 + 2^46 ) )   n = 46   d_n = 1+1i 
assign v[4'b0101] [46] = 21'h 0007FF;  // +1.9999999999999858 = 2^(47+1) *  1 * atan( 1 / (  1 + 2^47 ) )   n = 47   d_n = 1+1i 
assign v[4'b0101] [47] = 21'h 0007FF;  // +1.9999999999999929 = 2^(48+1) *  1 * atan( 1 / (  1 + 2^48 ) )   n = 48   d_n = 1+1i 
assign v[4'b0101] [48] = 21'h 0007FF;  // +1.9999999999999964 = 2^(49+1) *  1 * atan( 1 / (  1 + 2^49 ) )   n = 49   d_n = 1+1i 
assign v[4'b0101] [49] = 21'h 0007FF;  // +1.9999999999999982 = 2^(50+1) *  1 * atan( 1 / (  1 + 2^50 ) )   n = 50   d_n = 1+1i 
assign v[4'b0101] [50] = 21'h 0007FF;  // +1.9999999999999991 = 2^(51+1) *  1 * atan( 1 / (  1 + 2^51 ) )   n = 51   d_n = 1+1i 
assign v[4'b0101] [51] = 21'h 0007FF;  // +1.9999999999999996 = 2^(52+1) *  1 * atan( 1 / (  1 + 2^52 ) )   n = 52   d_n = 1+1i 
assign v[4'b0101] [52] = 21'h 000800;  // +2.0000000000000000 = 2^(53+1) *  1 * atan( 1 / (  1 + 2^53 ) )   n = 53   d_n = 1+1i 
assign v[4'b0101] [53] = 21'h 000800;  // +2.0000000000000000 = 2^(54+1) *  1 * atan( 1 / (  1 + 2^54 ) )   n = 54   d_n = 1+1i 
assign v[4'b0101] [54] = 21'h 000800;  // +2.0000000000000000 = 2^(55+1) *  1 * atan( 1 / (  1 + 2^55 ) )   n = 55   d_n = 1+1i 
assign v[4'b0101] [55] = 21'h 000800;  // +2.0000000000000000 = 2^(56+1) *  1 * atan( 1 / (  1 + 2^56 ) )   n = 56   d_n = 1+1i 
assign v[4'b0101] [56] = 21'h 000800;  // +2.0000000000000000 = 2^(57+1) *  1 * atan( 1 / (  1 + 2^57 ) )   n = 57   d_n = 1+1i 
assign v[4'b0101] [57] = 21'h 000800;  // +2.0000000000000000 = 2^(58+1) *  1 * atan( 1 / (  1 + 2^58 ) )   n = 58   d_n = 1+1i 
assign v[4'b0101] [58] = 21'h 000800;  // +2.0000000000000000 = 2^(59+1) *  1 * atan( 1 / (  1 + 2^59 ) )   n = 59   d_n = 1+1i 
assign v[4'b0101] [59] = 21'h 000800;  // +2.0000000000000000 = 2^(60+1) *  1 * atan( 1 / (  1 + 2^60 ) )   n = 60   d_n = 1+1i 
assign v[4'b0101] [60] = 21'h 000800;  // +2.0000000000000000 = 2^(61+1) *  1 * atan( 1 / (  1 + 2^61 ) )   n = 61   d_n = 1+1i 
assign v[4'b0101] [61] = 21'h 000800;  // +2.0000000000000000 = 2^(62+1) *  1 * atan( 1 / (  1 + 2^62 ) )   n = 62   d_n = 1+1i 
assign v[4'b0101] [62] = 21'h 000800;  // +2.0000000000000000 = 2^(63+1) *  1 * atan( 1 / (  1 + 2^63 ) )   n = 63   d_n = 1+1i 
assign v[4'b0101] [63] = 21'h 000800;  // +2.0000000000000000 = 2^(64+1) *  1 * atan( 1 / (  1 + 2^64 ) )   n = 64   d_n = 1+1i 
assign v[4'b0110] [00] = 21'h 00076B;  // +1.8545904360032244 = 2^(1+1) *  1 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = 0+1i 
assign v[4'b0110] [01] = 21'h 0007D6;  // +1.9598293050149131 = 2^(2+1) *  1 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = 0+1i 
assign v[4'b0110] [02] = 21'h 0007F5;  // +1.9896799127481830 = 2^(3+1) *  1 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = 0+1i 
assign v[4'b0110] [03] = 21'h 0007FD;  // +1.9974019198706352 = 2^(4+1) *  1 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = 0+1i 
assign v[4'b0110] [04] = 21'h 0007FF;  // +1.9993493395371698 = 2^(5+1) *  1 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = 0+1i 
assign v[4'b0110] [05] = 21'h 0007FF;  // +1.9998372634210344 = 2^(6+1) *  1 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = 0+1i 
assign v[4'b0110] [06] = 21'h 0007FF;  // +1.9999593113858845 = 2^(7+1) *  1 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = 0+1i 
assign v[4'b0110] [07] = 21'h 0007FF;  // +1.9999898275670895 = 2^(8+1) *  1 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = 0+1i 
assign v[4'b0110] [08] = 21'h 0007FF;  // +1.9999974568743104 = 2^(9+1) *  1 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = 0+1i 
assign v[4'b0110] [09] = 21'h 0007FF;  // +1.9999993642174863 = 2^(10+1) *  1 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = 0+1i 
assign v[4'b0110] [10] = 21'h 0007FF;  // +1.9999998410543034 = 2^(11+1) *  1 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = 0+1i 
assign v[4'b0110] [11] = 21'h 0007FF;  // +1.9999999602635716 = 2^(12+1) *  1 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = 0+1i 
assign v[4'b0110] [12] = 21'h 0007FF;  // +1.9999999900658927 = 2^(13+1) *  1 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = 0+1i 
assign v[4'b0110] [13] = 21'h 0007FF;  // +1.9999999975164731 = 2^(14+1) *  1 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = 0+1i 
assign v[4'b0110] [14] = 21'h 0007FF;  // +1.9999999993791182 = 2^(15+1) *  1 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = 0+1i 
assign v[4'b0110] [15] = 21'h 0007FF;  // +1.9999999998447795 = 2^(16+1) *  1 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = 0+1i 
assign v[4'b0110] [16] = 21'h 0007FF;  // +1.9999999999611948 = 2^(17+1) *  1 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = 0+1i 
assign v[4'b0110] [17] = 21'h 0007FF;  // +1.9999999999902986 = 2^(18+1) *  1 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = 0+1i 
assign v[4'b0110] [18] = 21'h 0007FF;  // +1.9999999999975746 = 2^(19+1) *  1 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = 0+1i 
assign v[4'b0110] [19] = 21'h 0007FF;  // +1.9999999999993936 = 2^(20+1) *  1 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = 0+1i 
assign v[4'b0110] [20] = 21'h 0007FF;  // +1.9999999999998483 = 2^(21+1) *  1 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = 0+1i 
assign v[4'b0110] [21] = 21'h 0007FF;  // +1.9999999999999620 = 2^(22+1) *  1 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = 0+1i 
assign v[4'b0110] [22] = 21'h 0007FF;  // +1.9999999999999905 = 2^(23+1) *  1 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = 0+1i 
assign v[4'b0110] [23] = 21'h 0007FF;  // +1.9999999999999976 = 2^(24+1) *  1 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = 0+1i 
assign v[4'b0110] [24] = 21'h 0007FF;  // +1.9999999999999993 = 2^(25+1) *  1 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = 0+1i 
assign v[4'b0110] [25] = 21'h 0007FF;  // +1.9999999999999998 = 2^(26+1) *  1 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = 0+1i 
assign v[4'b0110] [26] = 21'h 000800;  // +2.0000000000000000 = 2^(27+1) *  1 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = 0+1i 
assign v[4'b0110] [27] = 21'h 000800;  // +2.0000000000000000 = 2^(28+1) *  1 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = 0+1i 
assign v[4'b0110] [28] = 21'h 000800;  // +2.0000000000000000 = 2^(29+1) *  1 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = 0+1i 
assign v[4'b0110] [29] = 21'h 000800;  // +2.0000000000000000 = 2^(30+1) *  1 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = 0+1i 
assign v[4'b0110] [30] = 21'h 000800;  // +2.0000000000000000 = 2^(31+1) *  1 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = 0+1i 
assign v[4'b0110] [31] = 21'h 000800;  // +2.0000000000000000 = 2^(32+1) *  1 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = 0+1i 
assign v[4'b0110] [32] = 21'h 000800;  // +2.0000000000000000 = 2^(33+1) *  1 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = 0+1i 
assign v[4'b0110] [33] = 21'h 000800;  // +2.0000000000000000 = 2^(34+1) *  1 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = 0+1i 
assign v[4'b0110] [34] = 21'h 000800;  // +2.0000000000000000 = 2^(35+1) *  1 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = 0+1i 
assign v[4'b0110] [35] = 21'h 000800;  // +2.0000000000000000 = 2^(36+1) *  1 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = 0+1i 
assign v[4'b0110] [36] = 21'h 000800;  // +2.0000000000000000 = 2^(37+1) *  1 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = 0+1i 
assign v[4'b0110] [37] = 21'h 000800;  // +2.0000000000000000 = 2^(38+1) *  1 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = 0+1i 
assign v[4'b0110] [38] = 21'h 000800;  // +2.0000000000000000 = 2^(39+1) *  1 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = 0+1i 
assign v[4'b0110] [39] = 21'h 000800;  // +2.0000000000000000 = 2^(40+1) *  1 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = 0+1i 
assign v[4'b0110] [40] = 21'h 000800;  // +2.0000000000000000 = 2^(41+1) *  1 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = 0+1i 
assign v[4'b0110] [41] = 21'h 000800;  // +2.0000000000000000 = 2^(42+1) *  1 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = 0+1i 
assign v[4'b0110] [42] = 21'h 000800;  // +2.0000000000000000 = 2^(43+1) *  1 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = 0+1i 
assign v[4'b0110] [43] = 21'h 000800;  // +2.0000000000000000 = 2^(44+1) *  1 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = 0+1i 
assign v[4'b0110] [44] = 21'h 000800;  // +2.0000000000000000 = 2^(45+1) *  1 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = 0+1i 
assign v[4'b0110] [45] = 21'h 000800;  // +2.0000000000000000 = 2^(46+1) *  1 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = 0+1i 
assign v[4'b0110] [46] = 21'h 000800;  // +2.0000000000000000 = 2^(47+1) *  1 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = 0+1i 
assign v[4'b0110] [47] = 21'h 000800;  // +2.0000000000000000 = 2^(48+1) *  1 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = 0+1i 
assign v[4'b0110] [48] = 21'h 000800;  // +2.0000000000000000 = 2^(49+1) *  1 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = 0+1i 
assign v[4'b0110] [49] = 21'h 000800;  // +2.0000000000000000 = 2^(50+1) *  1 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = 0+1i 
assign v[4'b0110] [50] = 21'h 000800;  // +2.0000000000000000 = 2^(51+1) *  1 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = 0+1i 
assign v[4'b0110] [51] = 21'h 000800;  // +2.0000000000000000 = 2^(52+1) *  1 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = 0+1i 
assign v[4'b0110] [52] = 21'h 000800;  // +2.0000000000000000 = 2^(53+1) *  1 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = 0+1i 
assign v[4'b0110] [53] = 21'h 000800;  // +2.0000000000000000 = 2^(54+1) *  1 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = 0+1i 
assign v[4'b0110] [54] = 21'h 000800;  // +2.0000000000000000 = 2^(55+1) *  1 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = 0+1i 
assign v[4'b0110] [55] = 21'h 000800;  // +2.0000000000000000 = 2^(56+1) *  1 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = 0+1i 
assign v[4'b0110] [56] = 21'h 000800;  // +2.0000000000000000 = 2^(57+1) *  1 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = 0+1i 
assign v[4'b0110] [57] = 21'h 000800;  // +2.0000000000000000 = 2^(58+1) *  1 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = 0+1i 
assign v[4'b0110] [58] = 21'h 000800;  // +2.0000000000000000 = 2^(59+1) *  1 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = 0+1i 
assign v[4'b0110] [59] = 21'h 000800;  // +2.0000000000000000 = 2^(60+1) *  1 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = 0+1i 
assign v[4'b0110] [60] = 21'h 000800;  // +2.0000000000000000 = 2^(61+1) *  1 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = 0+1i 
assign v[4'b0110] [61] = 21'h 000800;  // +2.0000000000000000 = 2^(62+1) *  1 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = 0+1i 
assign v[4'b0110] [62] = 21'h 000800;  // +2.0000000000000000 = 2^(63+1) *  1 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = 0+1i 
assign v[4'b0110] [63] = 21'h 000800;  // +2.0000000000000000 = 2^(64+1) *  1 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = 0+1i 
assign v[4'b0111] [00] = 21'h 000C90;  // +3.1415926535897931 = 2^(1+1) *  1 * atan( 1 / ( -1 + 2^1 ) )   n =  1   d_n = -1+1i 
assign v[4'b0111] [01] = 21'h 000A4B;  // +2.5740044351731375 = 2^(2+1) *  1 * atan( 1 / ( -1 + 2^2 ) )   n =  2   d_n = -1+1i 
assign v[4'b0111] [02] = 21'h 000914;  // +2.2703528736666230 = 2^(3+1) *  1 * atan( 1 / ( -1 + 2^3 ) )   n =  3   d_n = -1+1i 
assign v[4'b0111] [03] = 21'h 000885;  // +2.1301812408263618 = 2^(4+1) *  1 * atan( 1 / ( -1 + 2^4 ) )   n =  4   d_n = -1+1i 
assign v[4'b0111] [04] = 21'h 000841;  // +2.0638004758562509 = 2^(5+1) *  1 * atan( 1 / ( -1 + 2^5 ) )   n =  5   d_n = -1+1i 
assign v[4'b0111] [05] = 21'h 000820;  // +2.0315754229491265 = 2^(6+1) *  1 * atan( 1 / ( -1 + 2^6 ) )   n =  6   d_n = -1+1i 
assign v[4'b0111] [06] = 21'h 000810;  // +2.0157063741697390 = 2^(7+1) *  1 * atan( 1 / ( -1 + 2^7 ) )   n =  7   d_n = -1+1i 
assign v[4'b0111] [07] = 21'h 000808;  // +2.0078328446771208 = 2^(8+1) *  1 * atan( 1 / ( -1 + 2^8 ) )   n =  8   d_n = -1+1i 
assign v[4'b0111] [08] = 21'h 000804;  // +2.0039113362396619 = 2^(9+1) *  1 * atan( 1 / ( -1 + 2^9 ) )   n =  9   d_n = -1+1i 
assign v[4'b0111] [09] = 21'h 000802;  // +2.0019543965642979 = 2^(10+1) *  1 * atan( 1 / ( -1 + 2^10 ) )   n = 10   d_n = -1+1i 
assign v[4'b0111] [10] = 21'h 000801;  // +2.0009768803913479 = 2^(11+1) *  1 * atan( 1 / ( -1 + 2^11 ) )   n = 11   d_n = -1+1i 
assign v[4'b0111] [11] = 21'h 000800;  // +2.0004883607228541 = 2^(12+1) *  1 * atan( 1 / ( -1 + 2^12 ) )   n = 12   d_n = -1+1i 
assign v[4'b0111] [12] = 21'h 000800;  // +2.0002441604932146 = 2^(13+1) *  1 * atan( 1 / ( -1 + 2^13 ) )   n = 13   d_n = -1+1i 
assign v[4'b0111] [13] = 21'h 000800;  // +2.0001220752795539 = 2^(14+1) *  1 * atan( 1 / ( -1 + 2^14 ) )   n = 14   d_n = -1+1i 
assign v[4'b0111] [14] = 21'h 000800;  // +2.0000610363980136 = 2^(15+1) *  1 * atan( 1 / ( -1 + 2^15 ) )   n = 15   d_n = -1+1i 
assign v[4'b0111] [15] = 21'h 000800;  // +2.0000305178885660 = 2^(16+1) *  1 * atan( 1 / ( -1 + 2^16 ) )   n = 16   d_n = -1+1i 
assign v[4'b0111] [16] = 21'h 000800;  // +2.0000152588666729 = 2^(17+1) *  1 * atan( 1 / ( -1 + 2^17 ) )   n = 17   d_n = -1+1i 
assign v[4'b0111] [17] = 21'h 000800;  // +2.0000076294139340 = 2^(18+1) *  1 * atan( 1 / ( -1 + 2^18 ) )   n = 18   d_n = -1+1i 
assign v[4'b0111] [18] = 21'h 000800;  // +2.0000038147021164 = 2^(19+1) *  1 * atan( 1 / ( -1 + 2^19 ) )   n = 19   d_n = -1+1i 
assign v[4'b0111] [19] = 21'h 000800;  // +2.0000019073498456 = 2^(20+1) *  1 * atan( 1 / ( -1 + 2^20 ) )   n = 20   d_n = -1+1i 
assign v[4'b0111] [20] = 21'h 000800;  // +2.0000009536746197 = 2^(21+1) *  1 * atan( 1 / ( -1 + 2^21 ) )   n = 21   d_n = -1+1i 
assign v[4'b0111] [21] = 21'h 000800;  // +2.0000004768372341 = 2^(22+1) *  1 * atan( 1 / ( -1 + 2^22 ) )   n = 22   d_n = -1+1i 
assign v[4'b0111] [22] = 21'h 000800;  // +2.0000002384185982 = 2^(23+1) *  1 * atan( 1 / ( -1 + 2^23 ) )   n = 23   d_n = -1+1i 
assign v[4'b0111] [23] = 21'h 000800;  // +2.0000001192092944 = 2^(24+1) *  1 * atan( 1 / ( -1 + 2^24 ) )   n = 24   d_n = -1+1i 
assign v[4'b0111] [24] = 21'h 000800;  // +2.0000000596046461 = 2^(25+1) *  1 * atan( 1 / ( -1 + 2^25 ) )   n = 25   d_n = -1+1i 
assign v[4'b0111] [25] = 21'h 000800;  // +2.0000000298023228 = 2^(26+1) *  1 * atan( 1 / ( -1 + 2^26 ) )   n = 26   d_n = -1+1i 
assign v[4'b0111] [26] = 21'h 000800;  // +2.0000000149011612 = 2^(27+1) *  1 * atan( 1 / ( -1 + 2^27 ) )   n = 27   d_n = -1+1i 
assign v[4'b0111] [27] = 21'h 000800;  // +2.0000000074505806 = 2^(28+1) *  1 * atan( 1 / ( -1 + 2^28 ) )   n = 28   d_n = -1+1i 
assign v[4'b0111] [28] = 21'h 000800;  // +2.0000000037252903 = 2^(29+1) *  1 * atan( 1 / ( -1 + 2^29 ) )   n = 29   d_n = -1+1i 
assign v[4'b0111] [29] = 21'h 000800;  // +2.0000000018626451 = 2^(30+1) *  1 * atan( 1 / ( -1 + 2^30 ) )   n = 30   d_n = -1+1i 
assign v[4'b0111] [30] = 21'h 000800;  // +2.0000000009313226 = 2^(31+1) *  1 * atan( 1 / ( -1 + 2^31 ) )   n = 31   d_n = -1+1i 
assign v[4'b0111] [31] = 21'h 000800;  // +2.0000000004656613 = 2^(32+1) *  1 * atan( 1 / ( -1 + 2^32 ) )   n = 32   d_n = -1+1i 
assign v[4'b0111] [32] = 21'h 000800;  // +2.0000000002328306 = 2^(33+1) *  1 * atan( 1 / ( -1 + 2^33 ) )   n = 33   d_n = -1+1i 
assign v[4'b0111] [33] = 21'h 000800;  // +2.0000000001164153 = 2^(34+1) *  1 * atan( 1 / ( -1 + 2^34 ) )   n = 34   d_n = -1+1i 
assign v[4'b0111] [34] = 21'h 000800;  // +2.0000000000582077 = 2^(35+1) *  1 * atan( 1 / ( -1 + 2^35 ) )   n = 35   d_n = -1+1i 
assign v[4'b0111] [35] = 21'h 000800;  // +2.0000000000291038 = 2^(36+1) *  1 * atan( 1 / ( -1 + 2^36 ) )   n = 36   d_n = -1+1i 
assign v[4'b0111] [36] = 21'h 000800;  // +2.0000000000145519 = 2^(37+1) *  1 * atan( 1 / ( -1 + 2^37 ) )   n = 37   d_n = -1+1i 
assign v[4'b0111] [37] = 21'h 000800;  // +2.0000000000072760 = 2^(38+1) *  1 * atan( 1 / ( -1 + 2^38 ) )   n = 38   d_n = -1+1i 
assign v[4'b0111] [38] = 21'h 000800;  // +2.0000000000036380 = 2^(39+1) *  1 * atan( 1 / ( -1 + 2^39 ) )   n = 39   d_n = -1+1i 
assign v[4'b0111] [39] = 21'h 000800;  // +2.0000000000018190 = 2^(40+1) *  1 * atan( 1 / ( -1 + 2^40 ) )   n = 40   d_n = -1+1i 
assign v[4'b0111] [40] = 21'h 000800;  // +2.0000000000009095 = 2^(41+1) *  1 * atan( 1 / ( -1 + 2^41 ) )   n = 41   d_n = -1+1i 
assign v[4'b0111] [41] = 21'h 000800;  // +2.0000000000004547 = 2^(42+1) *  1 * atan( 1 / ( -1 + 2^42 ) )   n = 42   d_n = -1+1i 
assign v[4'b0111] [42] = 21'h 000800;  // +2.0000000000002274 = 2^(43+1) *  1 * atan( 1 / ( -1 + 2^43 ) )   n = 43   d_n = -1+1i 
assign v[4'b0111] [43] = 21'h 000800;  // +2.0000000000001137 = 2^(44+1) *  1 * atan( 1 / ( -1 + 2^44 ) )   n = 44   d_n = -1+1i 
assign v[4'b0111] [44] = 21'h 000800;  // +2.0000000000000568 = 2^(45+1) *  1 * atan( 1 / ( -1 + 2^45 ) )   n = 45   d_n = -1+1i 
assign v[4'b0111] [45] = 21'h 000800;  // +2.0000000000000284 = 2^(46+1) *  1 * atan( 1 / ( -1 + 2^46 ) )   n = 46   d_n = -1+1i 
assign v[4'b0111] [46] = 21'h 000800;  // +2.0000000000000142 = 2^(47+1) *  1 * atan( 1 / ( -1 + 2^47 ) )   n = 47   d_n = -1+1i 
assign v[4'b0111] [47] = 21'h 000800;  // +2.0000000000000071 = 2^(48+1) *  1 * atan( 1 / ( -1 + 2^48 ) )   n = 48   d_n = -1+1i 
assign v[4'b0111] [48] = 21'h 000800;  // +2.0000000000000036 = 2^(49+1) *  1 * atan( 1 / ( -1 + 2^49 ) )   n = 49   d_n = -1+1i 
assign v[4'b0111] [49] = 21'h 000800;  // +2.0000000000000018 = 2^(50+1) *  1 * atan( 1 / ( -1 + 2^50 ) )   n = 50   d_n = -1+1i 
assign v[4'b0111] [50] = 21'h 000800;  // +2.0000000000000009 = 2^(51+1) *  1 * atan( 1 / ( -1 + 2^51 ) )   n = 51   d_n = -1+1i 
assign v[4'b0111] [51] = 21'h 000800;  // +2.0000000000000004 = 2^(52+1) *  1 * atan( 1 / ( -1 + 2^52 ) )   n = 52   d_n = -1+1i 
assign v[4'b0111] [52] = 21'h 000800;  // +2.0000000000000004 = 2^(53+1) *  1 * atan( 1 / ( -1 + 2^53 ) )   n = 53   d_n = -1+1i 
assign v[4'b0111] [53] = 21'h 000800;  // +2.0000000000000000 = 2^(54+1) *  1 * atan( 1 / ( -1 + 2^54 ) )   n = 54   d_n = -1+1i 
assign v[4'b0111] [54] = 21'h 000800;  // +2.0000000000000000 = 2^(55+1) *  1 * atan( 1 / ( -1 + 2^55 ) )   n = 55   d_n = -1+1i 
assign v[4'b0111] [55] = 21'h 000800;  // +2.0000000000000000 = 2^(56+1) *  1 * atan( 1 / ( -1 + 2^56 ) )   n = 56   d_n = -1+1i 
assign v[4'b0111] [56] = 21'h 000800;  // +2.0000000000000000 = 2^(57+1) *  1 * atan( 1 / ( -1 + 2^57 ) )   n = 57   d_n = -1+1i 
assign v[4'b0111] [57] = 21'h 000800;  // +2.0000000000000000 = 2^(58+1) *  1 * atan( 1 / ( -1 + 2^58 ) )   n = 58   d_n = -1+1i 
assign v[4'b0111] [58] = 21'h 000800;  // +2.0000000000000000 = 2^(59+1) *  1 * atan( 1 / ( -1 + 2^59 ) )   n = 59   d_n = -1+1i 
assign v[4'b0111] [59] = 21'h 000800;  // +2.0000000000000000 = 2^(60+1) *  1 * atan( 1 / ( -1 + 2^60 ) )   n = 60   d_n = -1+1i 
assign v[4'b0111] [60] = 21'h 000800;  // +2.0000000000000000 = 2^(61+1) *  1 * atan( 1 / ( -1 + 2^61 ) )   n = 61   d_n = -1+1i 
assign v[4'b0111] [61] = 21'h 000800;  // +2.0000000000000000 = 2^(62+1) *  1 * atan( 1 / ( -1 + 2^62 ) )   n = 62   d_n = -1+1i 
assign v[4'b0111] [62] = 21'h 000800;  // +2.0000000000000000 = 2^(63+1) *  1 * atan( 1 / ( -1 + 2^63 ) )   n = 63   d_n = -1+1i 
assign v[4'b0111] [63] = 21'h 000800;  // +2.0000000000000000 = 2^(64+1) *  1 * atan( 1 / ( -1 + 2^64 ) )   n = 64   d_n = -1+1i 
assign v[4'b1000] [00] = 21'h 000000;  // +0.0000000000000000 = 2^(1+1) *  0 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = 0 
assign v[4'b1000] [01] = 21'h 000000;  // +0.0000000000000000 = 2^(2+1) *  0 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = 0 
assign v[4'b1000] [02] = 21'h 000000;  // +0.0000000000000000 = 2^(3+1) *  0 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = 0 
assign v[4'b1000] [03] = 21'h 000000;  // +0.0000000000000000 = 2^(4+1) *  0 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = 0 
assign v[4'b1000] [04] = 21'h 000000;  // +0.0000000000000000 = 2^(5+1) *  0 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = 0 
assign v[4'b1000] [05] = 21'h 000000;  // +0.0000000000000000 = 2^(6+1) *  0 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = 0 
assign v[4'b1000] [06] = 21'h 000000;  // +0.0000000000000000 = 2^(7+1) *  0 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = 0 
assign v[4'b1000] [07] = 21'h 000000;  // +0.0000000000000000 = 2^(8+1) *  0 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = 0 
assign v[4'b1000] [08] = 21'h 000000;  // +0.0000000000000000 = 2^(9+1) *  0 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = 0 
assign v[4'b1000] [09] = 21'h 000000;  // +0.0000000000000000 = 2^(10+1) *  0 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = 0 
assign v[4'b1000] [10] = 21'h 000000;  // +0.0000000000000000 = 2^(11+1) *  0 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = 0 
assign v[4'b1000] [11] = 21'h 000000;  // +0.0000000000000000 = 2^(12+1) *  0 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = 0 
assign v[4'b1000] [12] = 21'h 000000;  // +0.0000000000000000 = 2^(13+1) *  0 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = 0 
assign v[4'b1000] [13] = 21'h 000000;  // +0.0000000000000000 = 2^(14+1) *  0 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = 0 
assign v[4'b1000] [14] = 21'h 000000;  // +0.0000000000000000 = 2^(15+1) *  0 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = 0 
assign v[4'b1000] [15] = 21'h 000000;  // +0.0000000000000000 = 2^(16+1) *  0 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = 0 
assign v[4'b1000] [16] = 21'h 000000;  // +0.0000000000000000 = 2^(17+1) *  0 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = 0 
assign v[4'b1000] [17] = 21'h 000000;  // +0.0000000000000000 = 2^(18+1) *  0 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = 0 
assign v[4'b1000] [18] = 21'h 000000;  // +0.0000000000000000 = 2^(19+1) *  0 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = 0 
assign v[4'b1000] [19] = 21'h 000000;  // +0.0000000000000000 = 2^(20+1) *  0 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = 0 
assign v[4'b1000] [20] = 21'h 000000;  // +0.0000000000000000 = 2^(21+1) *  0 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = 0 
assign v[4'b1000] [21] = 21'h 000000;  // +0.0000000000000000 = 2^(22+1) *  0 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = 0 
assign v[4'b1000] [22] = 21'h 000000;  // +0.0000000000000000 = 2^(23+1) *  0 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = 0 
assign v[4'b1000] [23] = 21'h 000000;  // +0.0000000000000000 = 2^(24+1) *  0 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = 0 
assign v[4'b1000] [24] = 21'h 000000;  // +0.0000000000000000 = 2^(25+1) *  0 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = 0 
assign v[4'b1000] [25] = 21'h 000000;  // +0.0000000000000000 = 2^(26+1) *  0 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = 0 
assign v[4'b1000] [26] = 21'h 000000;  // +0.0000000000000000 = 2^(27+1) *  0 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = 0 
assign v[4'b1000] [27] = 21'h 000000;  // +0.0000000000000000 = 2^(28+1) *  0 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = 0 
assign v[4'b1000] [28] = 21'h 000000;  // +0.0000000000000000 = 2^(29+1) *  0 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = 0 
assign v[4'b1000] [29] = 21'h 000000;  // +0.0000000000000000 = 2^(30+1) *  0 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = 0 
assign v[4'b1000] [30] = 21'h 000000;  // +0.0000000000000000 = 2^(31+1) *  0 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = 0 
assign v[4'b1000] [31] = 21'h 000000;  // +0.0000000000000000 = 2^(32+1) *  0 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = 0 
assign v[4'b1000] [32] = 21'h 000000;  // +0.0000000000000000 = 2^(33+1) *  0 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = 0 
assign v[4'b1000] [33] = 21'h 000000;  // +0.0000000000000000 = 2^(34+1) *  0 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = 0 
assign v[4'b1000] [34] = 21'h 000000;  // +0.0000000000000000 = 2^(35+1) *  0 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = 0 
assign v[4'b1000] [35] = 21'h 000000;  // +0.0000000000000000 = 2^(36+1) *  0 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = 0 
assign v[4'b1000] [36] = 21'h 000000;  // +0.0000000000000000 = 2^(37+1) *  0 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = 0 
assign v[4'b1000] [37] = 21'h 000000;  // +0.0000000000000000 = 2^(38+1) *  0 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = 0 
assign v[4'b1000] [38] = 21'h 000000;  // +0.0000000000000000 = 2^(39+1) *  0 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = 0 
assign v[4'b1000] [39] = 21'h 000000;  // +0.0000000000000000 = 2^(40+1) *  0 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = 0 
assign v[4'b1000] [40] = 21'h 000000;  // +0.0000000000000000 = 2^(41+1) *  0 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = 0 
assign v[4'b1000] [41] = 21'h 000000;  // +0.0000000000000000 = 2^(42+1) *  0 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = 0 
assign v[4'b1000] [42] = 21'h 000000;  // +0.0000000000000000 = 2^(43+1) *  0 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = 0 
assign v[4'b1000] [43] = 21'h 000000;  // +0.0000000000000000 = 2^(44+1) *  0 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = 0 
assign v[4'b1000] [44] = 21'h 000000;  // +0.0000000000000000 = 2^(45+1) *  0 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = 0 
assign v[4'b1000] [45] = 21'h 000000;  // +0.0000000000000000 = 2^(46+1) *  0 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = 0 
assign v[4'b1000] [46] = 21'h 000000;  // +0.0000000000000000 = 2^(47+1) *  0 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = 0 
assign v[4'b1000] [47] = 21'h 000000;  // +0.0000000000000000 = 2^(48+1) *  0 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = 0 
assign v[4'b1000] [48] = 21'h 000000;  // +0.0000000000000000 = 2^(49+1) *  0 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = 0 
assign v[4'b1000] [49] = 21'h 000000;  // +0.0000000000000000 = 2^(50+1) *  0 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = 0 
assign v[4'b1000] [50] = 21'h 000000;  // +0.0000000000000000 = 2^(51+1) *  0 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = 0 
assign v[4'b1000] [51] = 21'h 000000;  // +0.0000000000000000 = 2^(52+1) *  0 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = 0 
assign v[4'b1000] [52] = 21'h 000000;  // +0.0000000000000000 = 2^(53+1) *  0 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = 0 
assign v[4'b1000] [53] = 21'h 000000;  // +0.0000000000000000 = 2^(54+1) *  0 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = 0 
assign v[4'b1000] [54] = 21'h 000000;  // +0.0000000000000000 = 2^(55+1) *  0 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = 0 
assign v[4'b1000] [55] = 21'h 000000;  // +0.0000000000000000 = 2^(56+1) *  0 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = 0 
assign v[4'b1000] [56] = 21'h 000000;  // +0.0000000000000000 = 2^(57+1) *  0 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = 0 
assign v[4'b1000] [57] = 21'h 000000;  // +0.0000000000000000 = 2^(58+1) *  0 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = 0 
assign v[4'b1000] [58] = 21'h 000000;  // +0.0000000000000000 = 2^(59+1) *  0 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = 0 
assign v[4'b1000] [59] = 21'h 000000;  // +0.0000000000000000 = 2^(60+1) *  0 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = 0 
assign v[4'b1000] [60] = 21'h 000000;  // +0.0000000000000000 = 2^(61+1) *  0 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = 0 
assign v[4'b1000] [61] = 21'h 000000;  // +0.0000000000000000 = 2^(62+1) *  0 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = 0 
assign v[4'b1000] [62] = 21'h 000000;  // +0.0000000000000000 = 2^(63+1) *  0 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = 0 
assign v[4'b1000] [63] = 21'h 000000;  // +0.0000000000000000 = 2^(64+1) *  0 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = 0 
assign v[4'b1001] [00] = 21'h 000000;  // +0.0000000000000000 = 2^(1+1) *  0 * atan( 1 / (  1 + 2^1 ) )   n =  1   d_n = 1 
assign v[4'b1001] [01] = 21'h 000000;  // +0.0000000000000000 = 2^(2+1) *  0 * atan( 1 / (  1 + 2^2 ) )   n =  2   d_n = 1 
assign v[4'b1001] [02] = 21'h 000000;  // +0.0000000000000000 = 2^(3+1) *  0 * atan( 1 / (  1 + 2^3 ) )   n =  3   d_n = 1 
assign v[4'b1001] [03] = 21'h 000000;  // +0.0000000000000000 = 2^(4+1) *  0 * atan( 1 / (  1 + 2^4 ) )   n =  4   d_n = 1 
assign v[4'b1001] [04] = 21'h 000000;  // +0.0000000000000000 = 2^(5+1) *  0 * atan( 1 / (  1 + 2^5 ) )   n =  5   d_n = 1 
assign v[4'b1001] [05] = 21'h 000000;  // +0.0000000000000000 = 2^(6+1) *  0 * atan( 1 / (  1 + 2^6 ) )   n =  6   d_n = 1 
assign v[4'b1001] [06] = 21'h 000000;  // +0.0000000000000000 = 2^(7+1) *  0 * atan( 1 / (  1 + 2^7 ) )   n =  7   d_n = 1 
assign v[4'b1001] [07] = 21'h 000000;  // +0.0000000000000000 = 2^(8+1) *  0 * atan( 1 / (  1 + 2^8 ) )   n =  8   d_n = 1 
assign v[4'b1001] [08] = 21'h 000000;  // +0.0000000000000000 = 2^(9+1) *  0 * atan( 1 / (  1 + 2^9 ) )   n =  9   d_n = 1 
assign v[4'b1001] [09] = 21'h 000000;  // +0.0000000000000000 = 2^(10+1) *  0 * atan( 1 / (  1 + 2^10 ) )   n = 10   d_n = 1 
assign v[4'b1001] [10] = 21'h 000000;  // +0.0000000000000000 = 2^(11+1) *  0 * atan( 1 / (  1 + 2^11 ) )   n = 11   d_n = 1 
assign v[4'b1001] [11] = 21'h 000000;  // +0.0000000000000000 = 2^(12+1) *  0 * atan( 1 / (  1 + 2^12 ) )   n = 12   d_n = 1 
assign v[4'b1001] [12] = 21'h 000000;  // +0.0000000000000000 = 2^(13+1) *  0 * atan( 1 / (  1 + 2^13 ) )   n = 13   d_n = 1 
assign v[4'b1001] [13] = 21'h 000000;  // +0.0000000000000000 = 2^(14+1) *  0 * atan( 1 / (  1 + 2^14 ) )   n = 14   d_n = 1 
assign v[4'b1001] [14] = 21'h 000000;  // +0.0000000000000000 = 2^(15+1) *  0 * atan( 1 / (  1 + 2^15 ) )   n = 15   d_n = 1 
assign v[4'b1001] [15] = 21'h 000000;  // +0.0000000000000000 = 2^(16+1) *  0 * atan( 1 / (  1 + 2^16 ) )   n = 16   d_n = 1 
assign v[4'b1001] [16] = 21'h 000000;  // +0.0000000000000000 = 2^(17+1) *  0 * atan( 1 / (  1 + 2^17 ) )   n = 17   d_n = 1 
assign v[4'b1001] [17] = 21'h 000000;  // +0.0000000000000000 = 2^(18+1) *  0 * atan( 1 / (  1 + 2^18 ) )   n = 18   d_n = 1 
assign v[4'b1001] [18] = 21'h 000000;  // +0.0000000000000000 = 2^(19+1) *  0 * atan( 1 / (  1 + 2^19 ) )   n = 19   d_n = 1 
assign v[4'b1001] [19] = 21'h 000000;  // +0.0000000000000000 = 2^(20+1) *  0 * atan( 1 / (  1 + 2^20 ) )   n = 20   d_n = 1 
assign v[4'b1001] [20] = 21'h 000000;  // +0.0000000000000000 = 2^(21+1) *  0 * atan( 1 / (  1 + 2^21 ) )   n = 21   d_n = 1 
assign v[4'b1001] [21] = 21'h 000000;  // +0.0000000000000000 = 2^(22+1) *  0 * atan( 1 / (  1 + 2^22 ) )   n = 22   d_n = 1 
assign v[4'b1001] [22] = 21'h 000000;  // +0.0000000000000000 = 2^(23+1) *  0 * atan( 1 / (  1 + 2^23 ) )   n = 23   d_n = 1 
assign v[4'b1001] [23] = 21'h 000000;  // +0.0000000000000000 = 2^(24+1) *  0 * atan( 1 / (  1 + 2^24 ) )   n = 24   d_n = 1 
assign v[4'b1001] [24] = 21'h 000000;  // +0.0000000000000000 = 2^(25+1) *  0 * atan( 1 / (  1 + 2^25 ) )   n = 25   d_n = 1 
assign v[4'b1001] [25] = 21'h 000000;  // +0.0000000000000000 = 2^(26+1) *  0 * atan( 1 / (  1 + 2^26 ) )   n = 26   d_n = 1 
assign v[4'b1001] [26] = 21'h 000000;  // +0.0000000000000000 = 2^(27+1) *  0 * atan( 1 / (  1 + 2^27 ) )   n = 27   d_n = 1 
assign v[4'b1001] [27] = 21'h 000000;  // +0.0000000000000000 = 2^(28+1) *  0 * atan( 1 / (  1 + 2^28 ) )   n = 28   d_n = 1 
assign v[4'b1001] [28] = 21'h 000000;  // +0.0000000000000000 = 2^(29+1) *  0 * atan( 1 / (  1 + 2^29 ) )   n = 29   d_n = 1 
assign v[4'b1001] [29] = 21'h 000000;  // +0.0000000000000000 = 2^(30+1) *  0 * atan( 1 / (  1 + 2^30 ) )   n = 30   d_n = 1 
assign v[4'b1001] [30] = 21'h 000000;  // +0.0000000000000000 = 2^(31+1) *  0 * atan( 1 / (  1 + 2^31 ) )   n = 31   d_n = 1 
assign v[4'b1001] [31] = 21'h 000000;  // +0.0000000000000000 = 2^(32+1) *  0 * atan( 1 / (  1 + 2^32 ) )   n = 32   d_n = 1 
assign v[4'b1001] [32] = 21'h 000000;  // +0.0000000000000000 = 2^(33+1) *  0 * atan( 1 / (  1 + 2^33 ) )   n = 33   d_n = 1 
assign v[4'b1001] [33] = 21'h 000000;  // +0.0000000000000000 = 2^(34+1) *  0 * atan( 1 / (  1 + 2^34 ) )   n = 34   d_n = 1 
assign v[4'b1001] [34] = 21'h 000000;  // +0.0000000000000000 = 2^(35+1) *  0 * atan( 1 / (  1 + 2^35 ) )   n = 35   d_n = 1 
assign v[4'b1001] [35] = 21'h 000000;  // +0.0000000000000000 = 2^(36+1) *  0 * atan( 1 / (  1 + 2^36 ) )   n = 36   d_n = 1 
assign v[4'b1001] [36] = 21'h 000000;  // +0.0000000000000000 = 2^(37+1) *  0 * atan( 1 / (  1 + 2^37 ) )   n = 37   d_n = 1 
assign v[4'b1001] [37] = 21'h 000000;  // +0.0000000000000000 = 2^(38+1) *  0 * atan( 1 / (  1 + 2^38 ) )   n = 38   d_n = 1 
assign v[4'b1001] [38] = 21'h 000000;  // +0.0000000000000000 = 2^(39+1) *  0 * atan( 1 / (  1 + 2^39 ) )   n = 39   d_n = 1 
assign v[4'b1001] [39] = 21'h 000000;  // +0.0000000000000000 = 2^(40+1) *  0 * atan( 1 / (  1 + 2^40 ) )   n = 40   d_n = 1 
assign v[4'b1001] [40] = 21'h 000000;  // +0.0000000000000000 = 2^(41+1) *  0 * atan( 1 / (  1 + 2^41 ) )   n = 41   d_n = 1 
assign v[4'b1001] [41] = 21'h 000000;  // +0.0000000000000000 = 2^(42+1) *  0 * atan( 1 / (  1 + 2^42 ) )   n = 42   d_n = 1 
assign v[4'b1001] [42] = 21'h 000000;  // +0.0000000000000000 = 2^(43+1) *  0 * atan( 1 / (  1 + 2^43 ) )   n = 43   d_n = 1 
assign v[4'b1001] [43] = 21'h 000000;  // +0.0000000000000000 = 2^(44+1) *  0 * atan( 1 / (  1 + 2^44 ) )   n = 44   d_n = 1 
assign v[4'b1001] [44] = 21'h 000000;  // +0.0000000000000000 = 2^(45+1) *  0 * atan( 1 / (  1 + 2^45 ) )   n = 45   d_n = 1 
assign v[4'b1001] [45] = 21'h 000000;  // +0.0000000000000000 = 2^(46+1) *  0 * atan( 1 / (  1 + 2^46 ) )   n = 46   d_n = 1 
assign v[4'b1001] [46] = 21'h 000000;  // +0.0000000000000000 = 2^(47+1) *  0 * atan( 1 / (  1 + 2^47 ) )   n = 47   d_n = 1 
assign v[4'b1001] [47] = 21'h 000000;  // +0.0000000000000000 = 2^(48+1) *  0 * atan( 1 / (  1 + 2^48 ) )   n = 48   d_n = 1 
assign v[4'b1001] [48] = 21'h 000000;  // +0.0000000000000000 = 2^(49+1) *  0 * atan( 1 / (  1 + 2^49 ) )   n = 49   d_n = 1 
assign v[4'b1001] [49] = 21'h 000000;  // +0.0000000000000000 = 2^(50+1) *  0 * atan( 1 / (  1 + 2^50 ) )   n = 50   d_n = 1 
assign v[4'b1001] [50] = 21'h 000000;  // +0.0000000000000000 = 2^(51+1) *  0 * atan( 1 / (  1 + 2^51 ) )   n = 51   d_n = 1 
assign v[4'b1001] [51] = 21'h 000000;  // +0.0000000000000000 = 2^(52+1) *  0 * atan( 1 / (  1 + 2^52 ) )   n = 52   d_n = 1 
assign v[4'b1001] [52] = 21'h 000000;  // +0.0000000000000000 = 2^(53+1) *  0 * atan( 1 / (  1 + 2^53 ) )   n = 53   d_n = 1 
assign v[4'b1001] [53] = 21'h 000000;  // +0.0000000000000000 = 2^(54+1) *  0 * atan( 1 / (  1 + 2^54 ) )   n = 54   d_n = 1 
assign v[4'b1001] [54] = 21'h 000000;  // +0.0000000000000000 = 2^(55+1) *  0 * atan( 1 / (  1 + 2^55 ) )   n = 55   d_n = 1 
assign v[4'b1001] [55] = 21'h 000000;  // +0.0000000000000000 = 2^(56+1) *  0 * atan( 1 / (  1 + 2^56 ) )   n = 56   d_n = 1 
assign v[4'b1001] [56] = 21'h 000000;  // +0.0000000000000000 = 2^(57+1) *  0 * atan( 1 / (  1 + 2^57 ) )   n = 57   d_n = 1 
assign v[4'b1001] [57] = 21'h 000000;  // +0.0000000000000000 = 2^(58+1) *  0 * atan( 1 / (  1 + 2^58 ) )   n = 58   d_n = 1 
assign v[4'b1001] [58] = 21'h 000000;  // +0.0000000000000000 = 2^(59+1) *  0 * atan( 1 / (  1 + 2^59 ) )   n = 59   d_n = 1 
assign v[4'b1001] [59] = 21'h 000000;  // +0.0000000000000000 = 2^(60+1) *  0 * atan( 1 / (  1 + 2^60 ) )   n = 60   d_n = 1 
assign v[4'b1001] [60] = 21'h 000000;  // +0.0000000000000000 = 2^(61+1) *  0 * atan( 1 / (  1 + 2^61 ) )   n = 61   d_n = 1 
assign v[4'b1001] [61] = 21'h 000000;  // +0.0000000000000000 = 2^(62+1) *  0 * atan( 1 / (  1 + 2^62 ) )   n = 62   d_n = 1 
assign v[4'b1001] [62] = 21'h 000000;  // +0.0000000000000000 = 2^(63+1) *  0 * atan( 1 / (  1 + 2^63 ) )   n = 63   d_n = 1 
assign v[4'b1001] [63] = 21'h 000000;  // +0.0000000000000000 = 2^(64+1) *  0 * atan( 1 / (  1 + 2^64 ) )   n = 64   d_n = 1 
assign v[4'b1010] [00] = 21'h 000000;  // +0.0000000000000000 = 2^(1+1) *  0 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = -0 
assign v[4'b1010] [01] = 21'h 000000;  // +0.0000000000000000 = 2^(2+1) *  0 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = -0 
assign v[4'b1010] [02] = 21'h 000000;  // +0.0000000000000000 = 2^(3+1) *  0 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = -0 
assign v[4'b1010] [03] = 21'h 000000;  // +0.0000000000000000 = 2^(4+1) *  0 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = -0 
assign v[4'b1010] [04] = 21'h 000000;  // +0.0000000000000000 = 2^(5+1) *  0 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = -0 
assign v[4'b1010] [05] = 21'h 000000;  // +0.0000000000000000 = 2^(6+1) *  0 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = -0 
assign v[4'b1010] [06] = 21'h 000000;  // +0.0000000000000000 = 2^(7+1) *  0 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = -0 
assign v[4'b1010] [07] = 21'h 000000;  // +0.0000000000000000 = 2^(8+1) *  0 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = -0 
assign v[4'b1010] [08] = 21'h 000000;  // +0.0000000000000000 = 2^(9+1) *  0 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = -0 
assign v[4'b1010] [09] = 21'h 000000;  // +0.0000000000000000 = 2^(10+1) *  0 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = -0 
assign v[4'b1010] [10] = 21'h 000000;  // +0.0000000000000000 = 2^(11+1) *  0 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = -0 
assign v[4'b1010] [11] = 21'h 000000;  // +0.0000000000000000 = 2^(12+1) *  0 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = -0 
assign v[4'b1010] [12] = 21'h 000000;  // +0.0000000000000000 = 2^(13+1) *  0 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = -0 
assign v[4'b1010] [13] = 21'h 000000;  // +0.0000000000000000 = 2^(14+1) *  0 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = -0 
assign v[4'b1010] [14] = 21'h 000000;  // +0.0000000000000000 = 2^(15+1) *  0 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = -0 
assign v[4'b1010] [15] = 21'h 000000;  // +0.0000000000000000 = 2^(16+1) *  0 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = -0 
assign v[4'b1010] [16] = 21'h 000000;  // +0.0000000000000000 = 2^(17+1) *  0 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = -0 
assign v[4'b1010] [17] = 21'h 000000;  // +0.0000000000000000 = 2^(18+1) *  0 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = -0 
assign v[4'b1010] [18] = 21'h 000000;  // +0.0000000000000000 = 2^(19+1) *  0 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = -0 
assign v[4'b1010] [19] = 21'h 000000;  // +0.0000000000000000 = 2^(20+1) *  0 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = -0 
assign v[4'b1010] [20] = 21'h 000000;  // +0.0000000000000000 = 2^(21+1) *  0 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = -0 
assign v[4'b1010] [21] = 21'h 000000;  // +0.0000000000000000 = 2^(22+1) *  0 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = -0 
assign v[4'b1010] [22] = 21'h 000000;  // +0.0000000000000000 = 2^(23+1) *  0 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = -0 
assign v[4'b1010] [23] = 21'h 000000;  // +0.0000000000000000 = 2^(24+1) *  0 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = -0 
assign v[4'b1010] [24] = 21'h 000000;  // +0.0000000000000000 = 2^(25+1) *  0 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = -0 
assign v[4'b1010] [25] = 21'h 000000;  // +0.0000000000000000 = 2^(26+1) *  0 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = -0 
assign v[4'b1010] [26] = 21'h 000000;  // +0.0000000000000000 = 2^(27+1) *  0 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = -0 
assign v[4'b1010] [27] = 21'h 000000;  // +0.0000000000000000 = 2^(28+1) *  0 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = -0 
assign v[4'b1010] [28] = 21'h 000000;  // +0.0000000000000000 = 2^(29+1) *  0 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = -0 
assign v[4'b1010] [29] = 21'h 000000;  // +0.0000000000000000 = 2^(30+1) *  0 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = -0 
assign v[4'b1010] [30] = 21'h 000000;  // +0.0000000000000000 = 2^(31+1) *  0 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = -0 
assign v[4'b1010] [31] = 21'h 000000;  // +0.0000000000000000 = 2^(32+1) *  0 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = -0 
assign v[4'b1010] [32] = 21'h 000000;  // +0.0000000000000000 = 2^(33+1) *  0 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = -0 
assign v[4'b1010] [33] = 21'h 000000;  // +0.0000000000000000 = 2^(34+1) *  0 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = -0 
assign v[4'b1010] [34] = 21'h 000000;  // +0.0000000000000000 = 2^(35+1) *  0 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = -0 
assign v[4'b1010] [35] = 21'h 000000;  // +0.0000000000000000 = 2^(36+1) *  0 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = -0 
assign v[4'b1010] [36] = 21'h 000000;  // +0.0000000000000000 = 2^(37+1) *  0 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = -0 
assign v[4'b1010] [37] = 21'h 000000;  // +0.0000000000000000 = 2^(38+1) *  0 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = -0 
assign v[4'b1010] [38] = 21'h 000000;  // +0.0000000000000000 = 2^(39+1) *  0 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = -0 
assign v[4'b1010] [39] = 21'h 000000;  // +0.0000000000000000 = 2^(40+1) *  0 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = -0 
assign v[4'b1010] [40] = 21'h 000000;  // +0.0000000000000000 = 2^(41+1) *  0 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = -0 
assign v[4'b1010] [41] = 21'h 000000;  // +0.0000000000000000 = 2^(42+1) *  0 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = -0 
assign v[4'b1010] [42] = 21'h 000000;  // +0.0000000000000000 = 2^(43+1) *  0 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = -0 
assign v[4'b1010] [43] = 21'h 000000;  // +0.0000000000000000 = 2^(44+1) *  0 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = -0 
assign v[4'b1010] [44] = 21'h 000000;  // +0.0000000000000000 = 2^(45+1) *  0 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = -0 
assign v[4'b1010] [45] = 21'h 000000;  // +0.0000000000000000 = 2^(46+1) *  0 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = -0 
assign v[4'b1010] [46] = 21'h 000000;  // +0.0000000000000000 = 2^(47+1) *  0 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = -0 
assign v[4'b1010] [47] = 21'h 000000;  // +0.0000000000000000 = 2^(48+1) *  0 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = -0 
assign v[4'b1010] [48] = 21'h 000000;  // +0.0000000000000000 = 2^(49+1) *  0 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = -0 
assign v[4'b1010] [49] = 21'h 000000;  // +0.0000000000000000 = 2^(50+1) *  0 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = -0 
assign v[4'b1010] [50] = 21'h 000000;  // +0.0000000000000000 = 2^(51+1) *  0 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = -0 
assign v[4'b1010] [51] = 21'h 000000;  // +0.0000000000000000 = 2^(52+1) *  0 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = -0 
assign v[4'b1010] [52] = 21'h 000000;  // +0.0000000000000000 = 2^(53+1) *  0 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = -0 
assign v[4'b1010] [53] = 21'h 000000;  // +0.0000000000000000 = 2^(54+1) *  0 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = -0 
assign v[4'b1010] [54] = 21'h 000000;  // +0.0000000000000000 = 2^(55+1) *  0 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = -0 
assign v[4'b1010] [55] = 21'h 000000;  // +0.0000000000000000 = 2^(56+1) *  0 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = -0 
assign v[4'b1010] [56] = 21'h 000000;  // +0.0000000000000000 = 2^(57+1) *  0 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = -0 
assign v[4'b1010] [57] = 21'h 000000;  // +0.0000000000000000 = 2^(58+1) *  0 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = -0 
assign v[4'b1010] [58] = 21'h 000000;  // +0.0000000000000000 = 2^(59+1) *  0 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = -0 
assign v[4'b1010] [59] = 21'h 000000;  // +0.0000000000000000 = 2^(60+1) *  0 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = -0 
assign v[4'b1010] [60] = 21'h 000000;  // +0.0000000000000000 = 2^(61+1) *  0 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = -0 
assign v[4'b1010] [61] = 21'h 000000;  // +0.0000000000000000 = 2^(62+1) *  0 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = -0 
assign v[4'b1010] [62] = 21'h 000000;  // +0.0000000000000000 = 2^(63+1) *  0 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = -0 
assign v[4'b1010] [63] = 21'h 000000;  // +0.0000000000000000 = 2^(64+1) *  0 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = -0 
assign v[4'b1011] [00] = 21'h 000000;  // -0.0000000000000000 = 2^(1+1) *  0 * atan( 1 / ( -1 + 2^1 ) )   n =  1   d_n = -1 
assign v[4'b1011] [01] = 21'h 000000;  // -0.0000000000000000 = 2^(2+1) *  0 * atan( 1 / ( -1 + 2^2 ) )   n =  2   d_n = -1 
assign v[4'b1011] [02] = 21'h 000000;  // -0.0000000000000000 = 2^(3+1) *  0 * atan( 1 / ( -1 + 2^3 ) )   n =  3   d_n = -1 
assign v[4'b1011] [03] = 21'h 000000;  // -0.0000000000000000 = 2^(4+1) *  0 * atan( 1 / ( -1 + 2^4 ) )   n =  4   d_n = -1 
assign v[4'b1011] [04] = 21'h 000000;  // -0.0000000000000000 = 2^(5+1) *  0 * atan( 1 / ( -1 + 2^5 ) )   n =  5   d_n = -1 
assign v[4'b1011] [05] = 21'h 000000;  // -0.0000000000000000 = 2^(6+1) *  0 * atan( 1 / ( -1 + 2^6 ) )   n =  6   d_n = -1 
assign v[4'b1011] [06] = 21'h 000000;  // -0.0000000000000000 = 2^(7+1) *  0 * atan( 1 / ( -1 + 2^7 ) )   n =  7   d_n = -1 
assign v[4'b1011] [07] = 21'h 000000;  // -0.0000000000000000 = 2^(8+1) *  0 * atan( 1 / ( -1 + 2^8 ) )   n =  8   d_n = -1 
assign v[4'b1011] [08] = 21'h 000000;  // -0.0000000000000000 = 2^(9+1) *  0 * atan( 1 / ( -1 + 2^9 ) )   n =  9   d_n = -1 
assign v[4'b1011] [09] = 21'h 000000;  // -0.0000000000000000 = 2^(10+1) *  0 * atan( 1 / ( -1 + 2^10 ) )   n = 10   d_n = -1 
assign v[4'b1011] [10] = 21'h 000000;  // -0.0000000000000000 = 2^(11+1) *  0 * atan( 1 / ( -1 + 2^11 ) )   n = 11   d_n = -1 
assign v[4'b1011] [11] = 21'h 000000;  // -0.0000000000000000 = 2^(12+1) *  0 * atan( 1 / ( -1 + 2^12 ) )   n = 12   d_n = -1 
assign v[4'b1011] [12] = 21'h 000000;  // -0.0000000000000000 = 2^(13+1) *  0 * atan( 1 / ( -1 + 2^13 ) )   n = 13   d_n = -1 
assign v[4'b1011] [13] = 21'h 000000;  // -0.0000000000000000 = 2^(14+1) *  0 * atan( 1 / ( -1 + 2^14 ) )   n = 14   d_n = -1 
assign v[4'b1011] [14] = 21'h 000000;  // -0.0000000000000000 = 2^(15+1) *  0 * atan( 1 / ( -1 + 2^15 ) )   n = 15   d_n = -1 
assign v[4'b1011] [15] = 21'h 000000;  // -0.0000000000000000 = 2^(16+1) *  0 * atan( 1 / ( -1 + 2^16 ) )   n = 16   d_n = -1 
assign v[4'b1011] [16] = 21'h 000000;  // -0.0000000000000000 = 2^(17+1) *  0 * atan( 1 / ( -1 + 2^17 ) )   n = 17   d_n = -1 
assign v[4'b1011] [17] = 21'h 000000;  // -0.0000000000000000 = 2^(18+1) *  0 * atan( 1 / ( -1 + 2^18 ) )   n = 18   d_n = -1 
assign v[4'b1011] [18] = 21'h 000000;  // -0.0000000000000000 = 2^(19+1) *  0 * atan( 1 / ( -1 + 2^19 ) )   n = 19   d_n = -1 
assign v[4'b1011] [19] = 21'h 000000;  // -0.0000000000000000 = 2^(20+1) *  0 * atan( 1 / ( -1 + 2^20 ) )   n = 20   d_n = -1 
assign v[4'b1011] [20] = 21'h 000000;  // -0.0000000000000000 = 2^(21+1) *  0 * atan( 1 / ( -1 + 2^21 ) )   n = 21   d_n = -1 
assign v[4'b1011] [21] = 21'h 000000;  // -0.0000000000000000 = 2^(22+1) *  0 * atan( 1 / ( -1 + 2^22 ) )   n = 22   d_n = -1 
assign v[4'b1011] [22] = 21'h 000000;  // -0.0000000000000000 = 2^(23+1) *  0 * atan( 1 / ( -1 + 2^23 ) )   n = 23   d_n = -1 
assign v[4'b1011] [23] = 21'h 000000;  // -0.0000000000000000 = 2^(24+1) *  0 * atan( 1 / ( -1 + 2^24 ) )   n = 24   d_n = -1 
assign v[4'b1011] [24] = 21'h 000000;  // -0.0000000000000000 = 2^(25+1) *  0 * atan( 1 / ( -1 + 2^25 ) )   n = 25   d_n = -1 
assign v[4'b1011] [25] = 21'h 000000;  // -0.0000000000000000 = 2^(26+1) *  0 * atan( 1 / ( -1 + 2^26 ) )   n = 26   d_n = -1 
assign v[4'b1011] [26] = 21'h 000000;  // -0.0000000000000000 = 2^(27+1) *  0 * atan( 1 / ( -1 + 2^27 ) )   n = 27   d_n = -1 
assign v[4'b1011] [27] = 21'h 000000;  // -0.0000000000000000 = 2^(28+1) *  0 * atan( 1 / ( -1 + 2^28 ) )   n = 28   d_n = -1 
assign v[4'b1011] [28] = 21'h 000000;  // -0.0000000000000000 = 2^(29+1) *  0 * atan( 1 / ( -1 + 2^29 ) )   n = 29   d_n = -1 
assign v[4'b1011] [29] = 21'h 000000;  // -0.0000000000000000 = 2^(30+1) *  0 * atan( 1 / ( -1 + 2^30 ) )   n = 30   d_n = -1 
assign v[4'b1011] [30] = 21'h 000000;  // -0.0000000000000000 = 2^(31+1) *  0 * atan( 1 / ( -1 + 2^31 ) )   n = 31   d_n = -1 
assign v[4'b1011] [31] = 21'h 000000;  // -0.0000000000000000 = 2^(32+1) *  0 * atan( 1 / ( -1 + 2^32 ) )   n = 32   d_n = -1 
assign v[4'b1011] [32] = 21'h 000000;  // -0.0000000000000000 = 2^(33+1) *  0 * atan( 1 / ( -1 + 2^33 ) )   n = 33   d_n = -1 
assign v[4'b1011] [33] = 21'h 000000;  // -0.0000000000000000 = 2^(34+1) *  0 * atan( 1 / ( -1 + 2^34 ) )   n = 34   d_n = -1 
assign v[4'b1011] [34] = 21'h 000000;  // -0.0000000000000000 = 2^(35+1) *  0 * atan( 1 / ( -1 + 2^35 ) )   n = 35   d_n = -1 
assign v[4'b1011] [35] = 21'h 000000;  // -0.0000000000000000 = 2^(36+1) *  0 * atan( 1 / ( -1 + 2^36 ) )   n = 36   d_n = -1 
assign v[4'b1011] [36] = 21'h 000000;  // -0.0000000000000000 = 2^(37+1) *  0 * atan( 1 / ( -1 + 2^37 ) )   n = 37   d_n = -1 
assign v[4'b1011] [37] = 21'h 000000;  // -0.0000000000000000 = 2^(38+1) *  0 * atan( 1 / ( -1 + 2^38 ) )   n = 38   d_n = -1 
assign v[4'b1011] [38] = 21'h 000000;  // -0.0000000000000000 = 2^(39+1) *  0 * atan( 1 / ( -1 + 2^39 ) )   n = 39   d_n = -1 
assign v[4'b1011] [39] = 21'h 000000;  // -0.0000000000000000 = 2^(40+1) *  0 * atan( 1 / ( -1 + 2^40 ) )   n = 40   d_n = -1 
assign v[4'b1011] [40] = 21'h 000000;  // -0.0000000000000000 = 2^(41+1) *  0 * atan( 1 / ( -1 + 2^41 ) )   n = 41   d_n = -1 
assign v[4'b1011] [41] = 21'h 000000;  // -0.0000000000000000 = 2^(42+1) *  0 * atan( 1 / ( -1 + 2^42 ) )   n = 42   d_n = -1 
assign v[4'b1011] [42] = 21'h 000000;  // -0.0000000000000000 = 2^(43+1) *  0 * atan( 1 / ( -1 + 2^43 ) )   n = 43   d_n = -1 
assign v[4'b1011] [43] = 21'h 000000;  // -0.0000000000000000 = 2^(44+1) *  0 * atan( 1 / ( -1 + 2^44 ) )   n = 44   d_n = -1 
assign v[4'b1011] [44] = 21'h 000000;  // -0.0000000000000000 = 2^(45+1) *  0 * atan( 1 / ( -1 + 2^45 ) )   n = 45   d_n = -1 
assign v[4'b1011] [45] = 21'h 000000;  // -0.0000000000000000 = 2^(46+1) *  0 * atan( 1 / ( -1 + 2^46 ) )   n = 46   d_n = -1 
assign v[4'b1011] [46] = 21'h 000000;  // -0.0000000000000000 = 2^(47+1) *  0 * atan( 1 / ( -1 + 2^47 ) )   n = 47   d_n = -1 
assign v[4'b1011] [47] = 21'h 000000;  // -0.0000000000000000 = 2^(48+1) *  0 * atan( 1 / ( -1 + 2^48 ) )   n = 48   d_n = -1 
assign v[4'b1011] [48] = 21'h 000000;  // -0.0000000000000000 = 2^(49+1) *  0 * atan( 1 / ( -1 + 2^49 ) )   n = 49   d_n = -1 
assign v[4'b1011] [49] = 21'h 000000;  // -0.0000000000000000 = 2^(50+1) *  0 * atan( 1 / ( -1 + 2^50 ) )   n = 50   d_n = -1 
assign v[4'b1011] [50] = 21'h 000000;  // -0.0000000000000000 = 2^(51+1) *  0 * atan( 1 / ( -1 + 2^51 ) )   n = 51   d_n = -1 
assign v[4'b1011] [51] = 21'h 000000;  // -0.0000000000000000 = 2^(52+1) *  0 * atan( 1 / ( -1 + 2^52 ) )   n = 52   d_n = -1 
assign v[4'b1011] [52] = 21'h 000000;  // -0.0000000000000000 = 2^(53+1) *  0 * atan( 1 / ( -1 + 2^53 ) )   n = 53   d_n = -1 
assign v[4'b1011] [53] = 21'h 000000;  // -0.0000000000000000 = 2^(54+1) *  0 * atan( 1 / ( -1 + 2^54 ) )   n = 54   d_n = -1 
assign v[4'b1011] [54] = 21'h 000000;  // -0.0000000000000000 = 2^(55+1) *  0 * atan( 1 / ( -1 + 2^55 ) )   n = 55   d_n = -1 
assign v[4'b1011] [55] = 21'h 000000;  // -0.0000000000000000 = 2^(56+1) *  0 * atan( 1 / ( -1 + 2^56 ) )   n = 56   d_n = -1 
assign v[4'b1011] [56] = 21'h 000000;  // -0.0000000000000000 = 2^(57+1) *  0 * atan( 1 / ( -1 + 2^57 ) )   n = 57   d_n = -1 
assign v[4'b1011] [57] = 21'h 000000;  // -0.0000000000000000 = 2^(58+1) *  0 * atan( 1 / ( -1 + 2^58 ) )   n = 58   d_n = -1 
assign v[4'b1011] [58] = 21'h 000000;  // -0.0000000000000000 = 2^(59+1) *  0 * atan( 1 / ( -1 + 2^59 ) )   n = 59   d_n = -1 
assign v[4'b1011] [59] = 21'h 000000;  // -0.0000000000000000 = 2^(60+1) *  0 * atan( 1 / ( -1 + 2^60 ) )   n = 60   d_n = -1 
assign v[4'b1011] [60] = 21'h 000000;  // -0.0000000000000000 = 2^(61+1) *  0 * atan( 1 / ( -1 + 2^61 ) )   n = 61   d_n = -1 
assign v[4'b1011] [61] = 21'h 000000;  // -0.0000000000000000 = 2^(62+1) *  0 * atan( 1 / ( -1 + 2^62 ) )   n = 62   d_n = -1 
assign v[4'b1011] [62] = 21'h 000000;  // -0.0000000000000000 = 2^(63+1) *  0 * atan( 1 / ( -1 + 2^63 ) )   n = 63   d_n = -1 
assign v[4'b1011] [63] = 21'h 000000;  // -0.0000000000000000 = 2^(64+1) *  0 * atan( 1 / ( -1 + 2^64 ) )   n = 64   d_n = -1 
assign v[4'b1100] [00] = 21'h 1FF894;  // -1.8545904360032244 = 2^(1+1) * -1 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = -0-1i 
assign v[4'b1100] [01] = 21'h 1FF829;  // -1.9598293050149131 = 2^(2+1) * -1 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = -0-1i 
assign v[4'b1100] [02] = 21'h 1FF80A;  // -1.9896799127481830 = 2^(3+1) * -1 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = -0-1i 
assign v[4'b1100] [03] = 21'h 1FF802;  // -1.9974019198706352 = 2^(4+1) * -1 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = -0-1i 
assign v[4'b1100] [04] = 21'h 1FF800;  // -1.9993493395371698 = 2^(5+1) * -1 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = -0-1i 
assign v[4'b1100] [05] = 21'h 1FF800;  // -1.9998372634210344 = 2^(6+1) * -1 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = -0-1i 
assign v[4'b1100] [06] = 21'h 1FF800;  // -1.9999593113858845 = 2^(7+1) * -1 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = -0-1i 
assign v[4'b1100] [07] = 21'h 1FF800;  // -1.9999898275670895 = 2^(8+1) * -1 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = -0-1i 
assign v[4'b1100] [08] = 21'h 1FF800;  // -1.9999974568743104 = 2^(9+1) * -1 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = -0-1i 
assign v[4'b1100] [09] = 21'h 1FF800;  // -1.9999993642174863 = 2^(10+1) * -1 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = -0-1i 
assign v[4'b1100] [10] = 21'h 1FF800;  // -1.9999998410543034 = 2^(11+1) * -1 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = -0-1i 
assign v[4'b1100] [11] = 21'h 1FF800;  // -1.9999999602635716 = 2^(12+1) * -1 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = -0-1i 
assign v[4'b1100] [12] = 21'h 1FF800;  // -1.9999999900658927 = 2^(13+1) * -1 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = -0-1i 
assign v[4'b1100] [13] = 21'h 1FF800;  // -1.9999999975164731 = 2^(14+1) * -1 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = -0-1i 
assign v[4'b1100] [14] = 21'h 1FF800;  // -1.9999999993791182 = 2^(15+1) * -1 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = -0-1i 
assign v[4'b1100] [15] = 21'h 1FF800;  // -1.9999999998447795 = 2^(16+1) * -1 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = -0-1i 
assign v[4'b1100] [16] = 21'h 1FF800;  // -1.9999999999611948 = 2^(17+1) * -1 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = -0-1i 
assign v[4'b1100] [17] = 21'h 1FF800;  // -1.9999999999902986 = 2^(18+1) * -1 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = -0-1i 
assign v[4'b1100] [18] = 21'h 1FF800;  // -1.9999999999975746 = 2^(19+1) * -1 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = -0-1i 
assign v[4'b1100] [19] = 21'h 1FF800;  // -1.9999999999993936 = 2^(20+1) * -1 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = -0-1i 
assign v[4'b1100] [20] = 21'h 1FF800;  // -1.9999999999998483 = 2^(21+1) * -1 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = -0-1i 
assign v[4'b1100] [21] = 21'h 1FF800;  // -1.9999999999999620 = 2^(22+1) * -1 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = -0-1i 
assign v[4'b1100] [22] = 21'h 1FF800;  // -1.9999999999999905 = 2^(23+1) * -1 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = -0-1i 
assign v[4'b1100] [23] = 21'h 1FF800;  // -1.9999999999999976 = 2^(24+1) * -1 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = -0-1i 
assign v[4'b1100] [24] = 21'h 1FF800;  // -1.9999999999999993 = 2^(25+1) * -1 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = -0-1i 
assign v[4'b1100] [25] = 21'h 1FF800;  // -1.9999999999999998 = 2^(26+1) * -1 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = -0-1i 
assign v[4'b1100] [26] = 21'h 1FF800;  // -2.0000000000000000 = 2^(27+1) * -1 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = -0-1i 
assign v[4'b1100] [27] = 21'h 1FF800;  // -2.0000000000000000 = 2^(28+1) * -1 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = -0-1i 
assign v[4'b1100] [28] = 21'h 1FF800;  // -2.0000000000000000 = 2^(29+1) * -1 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = -0-1i 
assign v[4'b1100] [29] = 21'h 1FF800;  // -2.0000000000000000 = 2^(30+1) * -1 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = -0-1i 
assign v[4'b1100] [30] = 21'h 1FF800;  // -2.0000000000000000 = 2^(31+1) * -1 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = -0-1i 
assign v[4'b1100] [31] = 21'h 1FF800;  // -2.0000000000000000 = 2^(32+1) * -1 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = -0-1i 
assign v[4'b1100] [32] = 21'h 1FF800;  // -2.0000000000000000 = 2^(33+1) * -1 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = -0-1i 
assign v[4'b1100] [33] = 21'h 1FF800;  // -2.0000000000000000 = 2^(34+1) * -1 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = -0-1i 
assign v[4'b1100] [34] = 21'h 1FF800;  // -2.0000000000000000 = 2^(35+1) * -1 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = -0-1i 
assign v[4'b1100] [35] = 21'h 1FF800;  // -2.0000000000000000 = 2^(36+1) * -1 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = -0-1i 
assign v[4'b1100] [36] = 21'h 1FF800;  // -2.0000000000000000 = 2^(37+1) * -1 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = -0-1i 
assign v[4'b1100] [37] = 21'h 1FF800;  // -2.0000000000000000 = 2^(38+1) * -1 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = -0-1i 
assign v[4'b1100] [38] = 21'h 1FF800;  // -2.0000000000000000 = 2^(39+1) * -1 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = -0-1i 
assign v[4'b1100] [39] = 21'h 1FF800;  // -2.0000000000000000 = 2^(40+1) * -1 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = -0-1i 
assign v[4'b1100] [40] = 21'h 1FF800;  // -2.0000000000000000 = 2^(41+1) * -1 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = -0-1i 
assign v[4'b1100] [41] = 21'h 1FF800;  // -2.0000000000000000 = 2^(42+1) * -1 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = -0-1i 
assign v[4'b1100] [42] = 21'h 1FF800;  // -2.0000000000000000 = 2^(43+1) * -1 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = -0-1i 
assign v[4'b1100] [43] = 21'h 1FF800;  // -2.0000000000000000 = 2^(44+1) * -1 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = -0-1i 
assign v[4'b1100] [44] = 21'h 1FF800;  // -2.0000000000000000 = 2^(45+1) * -1 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = -0-1i 
assign v[4'b1100] [45] = 21'h 1FF800;  // -2.0000000000000000 = 2^(46+1) * -1 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = -0-1i 
assign v[4'b1100] [46] = 21'h 1FF800;  // -2.0000000000000000 = 2^(47+1) * -1 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = -0-1i 
assign v[4'b1100] [47] = 21'h 1FF800;  // -2.0000000000000000 = 2^(48+1) * -1 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = -0-1i 
assign v[4'b1100] [48] = 21'h 1FF800;  // -2.0000000000000000 = 2^(49+1) * -1 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = -0-1i 
assign v[4'b1100] [49] = 21'h 1FF800;  // -2.0000000000000000 = 2^(50+1) * -1 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = -0-1i 
assign v[4'b1100] [50] = 21'h 1FF800;  // -2.0000000000000000 = 2^(51+1) * -1 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = -0-1i 
assign v[4'b1100] [51] = 21'h 1FF800;  // -2.0000000000000000 = 2^(52+1) * -1 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = -0-1i 
assign v[4'b1100] [52] = 21'h 1FF800;  // -2.0000000000000000 = 2^(53+1) * -1 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = -0-1i 
assign v[4'b1100] [53] = 21'h 1FF800;  // -2.0000000000000000 = 2^(54+1) * -1 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = -0-1i 
assign v[4'b1100] [54] = 21'h 1FF800;  // -2.0000000000000000 = 2^(55+1) * -1 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = -0-1i 
assign v[4'b1100] [55] = 21'h 1FF800;  // -2.0000000000000000 = 2^(56+1) * -1 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = -0-1i 
assign v[4'b1100] [56] = 21'h 1FF800;  // -2.0000000000000000 = 2^(57+1) * -1 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = -0-1i 
assign v[4'b1100] [57] = 21'h 1FF800;  // -2.0000000000000000 = 2^(58+1) * -1 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = -0-1i 
assign v[4'b1100] [58] = 21'h 1FF800;  // -2.0000000000000000 = 2^(59+1) * -1 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = -0-1i 
assign v[4'b1100] [59] = 21'h 1FF800;  // -2.0000000000000000 = 2^(60+1) * -1 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = -0-1i 
assign v[4'b1100] [60] = 21'h 1FF800;  // -2.0000000000000000 = 2^(61+1) * -1 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = -0-1i 
assign v[4'b1100] [61] = 21'h 1FF800;  // -2.0000000000000000 = 2^(62+1) * -1 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = -0-1i 
assign v[4'b1100] [62] = 21'h 1FF800;  // -2.0000000000000000 = 2^(63+1) * -1 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = -0-1i 
assign v[4'b1100] [63] = 21'h 1FF800;  // -2.0000000000000000 = 2^(64+1) * -1 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = -0-1i 
assign v[4'b1101] [00] = 21'h 1FFADA;  // -1.2870022175865687 = 2^(1+1) * -1 * atan( 1 / (  1 + 2^1 ) )   n =  1   d_n = 1-1i 
assign v[4'b1101] [01] = 21'h 1FF9AE;  // -1.5791644787990460 = 2^(2+1) * -1 * atan( 1 / (  1 + 2^2 ) )   n =  2   d_n = 1-1i 
assign v[4'b1101] [02] = 21'h 1FF8EA;  // -1.7705155387823304 = 2^(3+1) * -1 * atan( 1 / (  1 + 2^3 ) )   n =  3   d_n = 1-1i 
assign v[4'b1101] [03] = 21'h 1FF87A;  // -1.8801863269031263 = 2^(4+1) * -1 * atan( 1 / (  1 + 2^4 ) )   n =  4   d_n = 1-1i 
assign v[4'b1101] [04] = 21'h 1FF83E;  // -1.9388006348016065 = 2^(5+1) * -1 * atan( 1 / (  1 + 2^5 ) )   n =  5   d_n = 1-1i 
assign v[4'b1101] [05] = 21'h 1FF81F;  // -1.9690754279161793 = 2^(6+1) * -1 * atan( 1 / (  1 + 2^6 ) )   n =  6   d_n = 1-1i 
assign v[4'b1101] [06] = 21'h 1FF80F;  // -1.9844563743249595 = 2^(7+1) * -1 * atan( 1 / (  1 + 2^7 ) )   n =  7   d_n = 1-1i 
assign v[4'b1101] [07] = 21'h 1FF807;  // -1.9922078446819715 = 2^(8+1) * -1 * atan( 1 / (  1 + 2^8 ) )   n =  8   d_n = 1-1i 
assign v[4'b1101] [08] = 21'h 1FF803;  // -1.9960988362398133 = 2^(9+1) * -1 * atan( 1 / (  1 + 2^9 ) )   n =  9   d_n = 1-1i 
assign v[4'b1101] [09] = 21'h 1FF801;  // -1.9980481465643023 = 2^(10+1) * -1 * atan( 1 / (  1 + 2^10 ) )   n = 10   d_n = 1-1i 
assign v[4'b1101] [10] = 21'h 1FF800;  // -1.9990237553913479 = 2^(11+1) * -1 * atan( 1 / (  1 + 2^11 ) )   n = 11   d_n = 1-1i 
assign v[4'b1101] [11] = 21'h 1FF800;  // -1.9995117982228541 = 2^(12+1) * -1 * atan( 1 / (  1 + 2^12 ) )   n = 12   d_n = 1-1i 
assign v[4'b1101] [12] = 21'h 1FF800;  // -1.9997558792432146 = 2^(13+1) * -1 * atan( 1 / (  1 + 2^13 ) )   n = 13   d_n = 1-1i 
assign v[4'b1101] [13] = 21'h 1FF800;  // -1.9998779346545537 = 2^(14+1) * -1 * atan( 1 / (  1 + 2^14 ) )   n = 14   d_n = 1-1i 
assign v[4'b1101] [14] = 21'h 1FF800;  // -1.9999389660855134 = 2^(15+1) * -1 * atan( 1 / (  1 + 2^15 ) )   n = 15   d_n = 1-1i 
assign v[4'b1101] [15] = 21'h 1FF800;  // -1.9999694827323158 = 2^(16+1) * -1 * atan( 1 / (  1 + 2^16 ) )   n = 16   d_n = 1-1i 
assign v[4'b1101] [16] = 21'h 1FF800;  // -1.9999847412885476 = 2^(17+1) * -1 * atan( 1 / (  1 + 2^17 ) )   n = 17   d_n = 1-1i 
assign v[4'b1101] [17] = 21'h 1FF800;  // -1.9999923706248712 = 2^(18+1) * -1 * atan( 1 / (  1 + 2^18 ) )   n = 18   d_n = 1-1i 
assign v[4'b1101] [18] = 21'h 1FF800;  // -1.9999961853075849 = 2^(19+1) * -1 * atan( 1 / (  1 + 2^19 ) )   n = 19   d_n = 1-1i 
assign v[4'b1101] [19] = 21'h 1FF800;  // -1.9999980926525798 = 2^(20+1) * -1 * atan( 1 / (  1 + 2^20 ) )   n = 20   d_n = 1-1i 
assign v[4'b1101] [20] = 21'h 1FF800;  // -1.9999990463259867 = 2^(21+1) * -1 * atan( 1 / (  1 + 2^21 ) )   n = 21   d_n = 1-1i 
assign v[4'b1101] [21] = 21'h 1FF800;  // -1.9999995231629175 = 2^(22+1) * -1 * atan( 1 / (  1 + 2^22 ) )   n = 22   d_n = 1-1i 
assign v[4'b1101] [22] = 21'h 1FF800;  // -1.9999997615814398 = 2^(23+1) * -1 * atan( 1 / (  1 + 2^23 ) )   n = 23   d_n = 1-1i 
assign v[4'b1101] [23] = 21'h 1FF800;  // -1.9999998807907151 = 2^(24+1) * -1 * atan( 1 / (  1 + 2^24 ) )   n = 24   d_n = 1-1i 
assign v[4'b1101] [24] = 21'h 1FF800;  // -1.9999999403953563 = 2^(25+1) * -1 * atan( 1 / (  1 + 2^25 ) )   n = 25   d_n = 1-1i 
assign v[4'b1101] [25] = 21'h 1FF800;  // -1.9999999701976778 = 2^(26+1) * -1 * atan( 1 / (  1 + 2^26 ) )   n = 26   d_n = 1-1i 
assign v[4'b1101] [26] = 21'h 1FF800;  // -1.9999999850988388 = 2^(27+1) * -1 * atan( 1 / (  1 + 2^27 ) )   n = 27   d_n = 1-1i 
assign v[4'b1101] [27] = 21'h 1FF800;  // -1.9999999925494194 = 2^(28+1) * -1 * atan( 1 / (  1 + 2^28 ) )   n = 28   d_n = 1-1i 
assign v[4'b1101] [28] = 21'h 1FF800;  // -1.9999999962747097 = 2^(29+1) * -1 * atan( 1 / (  1 + 2^29 ) )   n = 29   d_n = 1-1i 
assign v[4'b1101] [29] = 21'h 1FF800;  // -1.9999999981373549 = 2^(30+1) * -1 * atan( 1 / (  1 + 2^30 ) )   n = 30   d_n = 1-1i 
assign v[4'b1101] [30] = 21'h 1FF800;  // -1.9999999990686774 = 2^(31+1) * -1 * atan( 1 / (  1 + 2^31 ) )   n = 31   d_n = 1-1i 
assign v[4'b1101] [31] = 21'h 1FF800;  // -1.9999999995343387 = 2^(32+1) * -1 * atan( 1 / (  1 + 2^32 ) )   n = 32   d_n = 1-1i 
assign v[4'b1101] [32] = 21'h 1FF800;  // -1.9999999997671694 = 2^(33+1) * -1 * atan( 1 / (  1 + 2^33 ) )   n = 33   d_n = 1-1i 
assign v[4'b1101] [33] = 21'h 1FF800;  // -1.9999999998835847 = 2^(34+1) * -1 * atan( 1 / (  1 + 2^34 ) )   n = 34   d_n = 1-1i 
assign v[4'b1101] [34] = 21'h 1FF800;  // -1.9999999999417923 = 2^(35+1) * -1 * atan( 1 / (  1 + 2^35 ) )   n = 35   d_n = 1-1i 
assign v[4'b1101] [35] = 21'h 1FF800;  // -1.9999999999708962 = 2^(36+1) * -1 * atan( 1 / (  1 + 2^36 ) )   n = 36   d_n = 1-1i 
assign v[4'b1101] [36] = 21'h 1FF800;  // -1.9999999999854481 = 2^(37+1) * -1 * atan( 1 / (  1 + 2^37 ) )   n = 37   d_n = 1-1i 
assign v[4'b1101] [37] = 21'h 1FF800;  // -1.9999999999927240 = 2^(38+1) * -1 * atan( 1 / (  1 + 2^38 ) )   n = 38   d_n = 1-1i 
assign v[4'b1101] [38] = 21'h 1FF800;  // -1.9999999999963620 = 2^(39+1) * -1 * atan( 1 / (  1 + 2^39 ) )   n = 39   d_n = 1-1i 
assign v[4'b1101] [39] = 21'h 1FF800;  // -1.9999999999981810 = 2^(40+1) * -1 * atan( 1 / (  1 + 2^40 ) )   n = 40   d_n = 1-1i 
assign v[4'b1101] [40] = 21'h 1FF800;  // -1.9999999999990905 = 2^(41+1) * -1 * atan( 1 / (  1 + 2^41 ) )   n = 41   d_n = 1-1i 
assign v[4'b1101] [41] = 21'h 1FF800;  // -1.9999999999995453 = 2^(42+1) * -1 * atan( 1 / (  1 + 2^42 ) )   n = 42   d_n = 1-1i 
assign v[4'b1101] [42] = 21'h 1FF800;  // -1.9999999999997726 = 2^(43+1) * -1 * atan( 1 / (  1 + 2^43 ) )   n = 43   d_n = 1-1i 
assign v[4'b1101] [43] = 21'h 1FF800;  // -1.9999999999998863 = 2^(44+1) * -1 * atan( 1 / (  1 + 2^44 ) )   n = 44   d_n = 1-1i 
assign v[4'b1101] [44] = 21'h 1FF800;  // -1.9999999999999432 = 2^(45+1) * -1 * atan( 1 / (  1 + 2^45 ) )   n = 45   d_n = 1-1i 
assign v[4'b1101] [45] = 21'h 1FF800;  // -1.9999999999999716 = 2^(46+1) * -1 * atan( 1 / (  1 + 2^46 ) )   n = 46   d_n = 1-1i 
assign v[4'b1101] [46] = 21'h 1FF800;  // -1.9999999999999858 = 2^(47+1) * -1 * atan( 1 / (  1 + 2^47 ) )   n = 47   d_n = 1-1i 
assign v[4'b1101] [47] = 21'h 1FF800;  // -1.9999999999999929 = 2^(48+1) * -1 * atan( 1 / (  1 + 2^48 ) )   n = 48   d_n = 1-1i 
assign v[4'b1101] [48] = 21'h 1FF800;  // -1.9999999999999964 = 2^(49+1) * -1 * atan( 1 / (  1 + 2^49 ) )   n = 49   d_n = 1-1i 
assign v[4'b1101] [49] = 21'h 1FF800;  // -1.9999999999999982 = 2^(50+1) * -1 * atan( 1 / (  1 + 2^50 ) )   n = 50   d_n = 1-1i 
assign v[4'b1101] [50] = 21'h 1FF800;  // -1.9999999999999991 = 2^(51+1) * -1 * atan( 1 / (  1 + 2^51 ) )   n = 51   d_n = 1-1i 
assign v[4'b1101] [51] = 21'h 1FF800;  // -1.9999999999999996 = 2^(52+1) * -1 * atan( 1 / (  1 + 2^52 ) )   n = 52   d_n = 1-1i 
assign v[4'b1101] [52] = 21'h 1FF800;  // -2.0000000000000000 = 2^(53+1) * -1 * atan( 1 / (  1 + 2^53 ) )   n = 53   d_n = 1-1i 
assign v[4'b1101] [53] = 21'h 1FF800;  // -2.0000000000000000 = 2^(54+1) * -1 * atan( 1 / (  1 + 2^54 ) )   n = 54   d_n = 1-1i 
assign v[4'b1101] [54] = 21'h 1FF800;  // -2.0000000000000000 = 2^(55+1) * -1 * atan( 1 / (  1 + 2^55 ) )   n = 55   d_n = 1-1i 
assign v[4'b1101] [55] = 21'h 1FF800;  // -2.0000000000000000 = 2^(56+1) * -1 * atan( 1 / (  1 + 2^56 ) )   n = 56   d_n = 1-1i 
assign v[4'b1101] [56] = 21'h 1FF800;  // -2.0000000000000000 = 2^(57+1) * -1 * atan( 1 / (  1 + 2^57 ) )   n = 57   d_n = 1-1i 
assign v[4'b1101] [57] = 21'h 1FF800;  // -2.0000000000000000 = 2^(58+1) * -1 * atan( 1 / (  1 + 2^58 ) )   n = 58   d_n = 1-1i 
assign v[4'b1101] [58] = 21'h 1FF800;  // -2.0000000000000000 = 2^(59+1) * -1 * atan( 1 / (  1 + 2^59 ) )   n = 59   d_n = 1-1i 
assign v[4'b1101] [59] = 21'h 1FF800;  // -2.0000000000000000 = 2^(60+1) * -1 * atan( 1 / (  1 + 2^60 ) )   n = 60   d_n = 1-1i 
assign v[4'b1101] [60] = 21'h 1FF800;  // -2.0000000000000000 = 2^(61+1) * -1 * atan( 1 / (  1 + 2^61 ) )   n = 61   d_n = 1-1i 
assign v[4'b1101] [61] = 21'h 1FF800;  // -2.0000000000000000 = 2^(62+1) * -1 * atan( 1 / (  1 + 2^62 ) )   n = 62   d_n = 1-1i 
assign v[4'b1101] [62] = 21'h 1FF800;  // -2.0000000000000000 = 2^(63+1) * -1 * atan( 1 / (  1 + 2^63 ) )   n = 63   d_n = 1-1i 
assign v[4'b1101] [63] = 21'h 1FF800;  // -2.0000000000000000 = 2^(64+1) * -1 * atan( 1 / (  1 + 2^64 ) )   n = 64   d_n = 1-1i 
assign v[4'b1110] [00] = 21'h 1FF894;  // -1.8545904360032244 = 2^(1+1) * -1 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = -0-1i 
assign v[4'b1110] [01] = 21'h 1FF829;  // -1.9598293050149131 = 2^(2+1) * -1 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = -0-1i 
assign v[4'b1110] [02] = 21'h 1FF80A;  // -1.9896799127481830 = 2^(3+1) * -1 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = -0-1i 
assign v[4'b1110] [03] = 21'h 1FF802;  // -1.9974019198706352 = 2^(4+1) * -1 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = -0-1i 
assign v[4'b1110] [04] = 21'h 1FF800;  // -1.9993493395371698 = 2^(5+1) * -1 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = -0-1i 
assign v[4'b1110] [05] = 21'h 1FF800;  // -1.9998372634210344 = 2^(6+1) * -1 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = -0-1i 
assign v[4'b1110] [06] = 21'h 1FF800;  // -1.9999593113858845 = 2^(7+1) * -1 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = -0-1i 
assign v[4'b1110] [07] = 21'h 1FF800;  // -1.9999898275670895 = 2^(8+1) * -1 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = -0-1i 
assign v[4'b1110] [08] = 21'h 1FF800;  // -1.9999974568743104 = 2^(9+1) * -1 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = -0-1i 
assign v[4'b1110] [09] = 21'h 1FF800;  // -1.9999993642174863 = 2^(10+1) * -1 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = -0-1i 
assign v[4'b1110] [10] = 21'h 1FF800;  // -1.9999998410543034 = 2^(11+1) * -1 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = -0-1i 
assign v[4'b1110] [11] = 21'h 1FF800;  // -1.9999999602635716 = 2^(12+1) * -1 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = -0-1i 
assign v[4'b1110] [12] = 21'h 1FF800;  // -1.9999999900658927 = 2^(13+1) * -1 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = -0-1i 
assign v[4'b1110] [13] = 21'h 1FF800;  // -1.9999999975164731 = 2^(14+1) * -1 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = -0-1i 
assign v[4'b1110] [14] = 21'h 1FF800;  // -1.9999999993791182 = 2^(15+1) * -1 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = -0-1i 
assign v[4'b1110] [15] = 21'h 1FF800;  // -1.9999999998447795 = 2^(16+1) * -1 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = -0-1i 
assign v[4'b1110] [16] = 21'h 1FF800;  // -1.9999999999611948 = 2^(17+1) * -1 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = -0-1i 
assign v[4'b1110] [17] = 21'h 1FF800;  // -1.9999999999902986 = 2^(18+1) * -1 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = -0-1i 
assign v[4'b1110] [18] = 21'h 1FF800;  // -1.9999999999975746 = 2^(19+1) * -1 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = -0-1i 
assign v[4'b1110] [19] = 21'h 1FF800;  // -1.9999999999993936 = 2^(20+1) * -1 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = -0-1i 
assign v[4'b1110] [20] = 21'h 1FF800;  // -1.9999999999998483 = 2^(21+1) * -1 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = -0-1i 
assign v[4'b1110] [21] = 21'h 1FF800;  // -1.9999999999999620 = 2^(22+1) * -1 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = -0-1i 
assign v[4'b1110] [22] = 21'h 1FF800;  // -1.9999999999999905 = 2^(23+1) * -1 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = -0-1i 
assign v[4'b1110] [23] = 21'h 1FF800;  // -1.9999999999999976 = 2^(24+1) * -1 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = -0-1i 
assign v[4'b1110] [24] = 21'h 1FF800;  // -1.9999999999999993 = 2^(25+1) * -1 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = -0-1i 
assign v[4'b1110] [25] = 21'h 1FF800;  // -1.9999999999999998 = 2^(26+1) * -1 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = -0-1i 
assign v[4'b1110] [26] = 21'h 1FF800;  // -2.0000000000000000 = 2^(27+1) * -1 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = -0-1i 
assign v[4'b1110] [27] = 21'h 1FF800;  // -2.0000000000000000 = 2^(28+1) * -1 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = -0-1i 
assign v[4'b1110] [28] = 21'h 1FF800;  // -2.0000000000000000 = 2^(29+1) * -1 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = -0-1i 
assign v[4'b1110] [29] = 21'h 1FF800;  // -2.0000000000000000 = 2^(30+1) * -1 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = -0-1i 
assign v[4'b1110] [30] = 21'h 1FF800;  // -2.0000000000000000 = 2^(31+1) * -1 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = -0-1i 
assign v[4'b1110] [31] = 21'h 1FF800;  // -2.0000000000000000 = 2^(32+1) * -1 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = -0-1i 
assign v[4'b1110] [32] = 21'h 1FF800;  // -2.0000000000000000 = 2^(33+1) * -1 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = -0-1i 
assign v[4'b1110] [33] = 21'h 1FF800;  // -2.0000000000000000 = 2^(34+1) * -1 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = -0-1i 
assign v[4'b1110] [34] = 21'h 1FF800;  // -2.0000000000000000 = 2^(35+1) * -1 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = -0-1i 
assign v[4'b1110] [35] = 21'h 1FF800;  // -2.0000000000000000 = 2^(36+1) * -1 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = -0-1i 
assign v[4'b1110] [36] = 21'h 1FF800;  // -2.0000000000000000 = 2^(37+1) * -1 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = -0-1i 
assign v[4'b1110] [37] = 21'h 1FF800;  // -2.0000000000000000 = 2^(38+1) * -1 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = -0-1i 
assign v[4'b1110] [38] = 21'h 1FF800;  // -2.0000000000000000 = 2^(39+1) * -1 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = -0-1i 
assign v[4'b1110] [39] = 21'h 1FF800;  // -2.0000000000000000 = 2^(40+1) * -1 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = -0-1i 
assign v[4'b1110] [40] = 21'h 1FF800;  // -2.0000000000000000 = 2^(41+1) * -1 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = -0-1i 
assign v[4'b1110] [41] = 21'h 1FF800;  // -2.0000000000000000 = 2^(42+1) * -1 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = -0-1i 
assign v[4'b1110] [42] = 21'h 1FF800;  // -2.0000000000000000 = 2^(43+1) * -1 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = -0-1i 
assign v[4'b1110] [43] = 21'h 1FF800;  // -2.0000000000000000 = 2^(44+1) * -1 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = -0-1i 
assign v[4'b1110] [44] = 21'h 1FF800;  // -2.0000000000000000 = 2^(45+1) * -1 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = -0-1i 
assign v[4'b1110] [45] = 21'h 1FF800;  // -2.0000000000000000 = 2^(46+1) * -1 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = -0-1i 
assign v[4'b1110] [46] = 21'h 1FF800;  // -2.0000000000000000 = 2^(47+1) * -1 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = -0-1i 
assign v[4'b1110] [47] = 21'h 1FF800;  // -2.0000000000000000 = 2^(48+1) * -1 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = -0-1i 
assign v[4'b1110] [48] = 21'h 1FF800;  // -2.0000000000000000 = 2^(49+1) * -1 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = -0-1i 
assign v[4'b1110] [49] = 21'h 1FF800;  // -2.0000000000000000 = 2^(50+1) * -1 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = -0-1i 
assign v[4'b1110] [50] = 21'h 1FF800;  // -2.0000000000000000 = 2^(51+1) * -1 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = -0-1i 
assign v[4'b1110] [51] = 21'h 1FF800;  // -2.0000000000000000 = 2^(52+1) * -1 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = -0-1i 
assign v[4'b1110] [52] = 21'h 1FF800;  // -2.0000000000000000 = 2^(53+1) * -1 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = -0-1i 
assign v[4'b1110] [53] = 21'h 1FF800;  // -2.0000000000000000 = 2^(54+1) * -1 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = -0-1i 
assign v[4'b1110] [54] = 21'h 1FF800;  // -2.0000000000000000 = 2^(55+1) * -1 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = -0-1i 
assign v[4'b1110] [55] = 21'h 1FF800;  // -2.0000000000000000 = 2^(56+1) * -1 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = -0-1i 
assign v[4'b1110] [56] = 21'h 1FF800;  // -2.0000000000000000 = 2^(57+1) * -1 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = -0-1i 
assign v[4'b1110] [57] = 21'h 1FF800;  // -2.0000000000000000 = 2^(58+1) * -1 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = -0-1i 
assign v[4'b1110] [58] = 21'h 1FF800;  // -2.0000000000000000 = 2^(59+1) * -1 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = -0-1i 
assign v[4'b1110] [59] = 21'h 1FF800;  // -2.0000000000000000 = 2^(60+1) * -1 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = -0-1i 
assign v[4'b1110] [60] = 21'h 1FF800;  // -2.0000000000000000 = 2^(61+1) * -1 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = -0-1i 
assign v[4'b1110] [61] = 21'h 1FF800;  // -2.0000000000000000 = 2^(62+1) * -1 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = -0-1i 
assign v[4'b1110] [62] = 21'h 1FF800;  // -2.0000000000000000 = 2^(63+1) * -1 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = -0-1i 
assign v[4'b1110] [63] = 21'h 1FF800;  // -2.0000000000000000 = 2^(64+1) * -1 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = -0-1i 
assign v[4'b1111] [00] = 21'h 1FF36F;  // -3.1415926535897931 = 2^(1+1) * -1 * atan( 1 / ( -1 + 2^1 ) )   n =  1   d_n = -1-1i 
assign v[4'b1111] [01] = 21'h 1FF5B4;  // -2.5740044351731375 = 2^(2+1) * -1 * atan( 1 / ( -1 + 2^2 ) )   n =  2   d_n = -1-1i 
assign v[4'b1111] [02] = 21'h 1FF6EB;  // -2.2703528736666230 = 2^(3+1) * -1 * atan( 1 / ( -1 + 2^3 ) )   n =  3   d_n = -1-1i 
assign v[4'b1111] [03] = 21'h 1FF77A;  // -2.1301812408263618 = 2^(4+1) * -1 * atan( 1 / ( -1 + 2^4 ) )   n =  4   d_n = -1-1i 
assign v[4'b1111] [04] = 21'h 1FF7BE;  // -2.0638004758562509 = 2^(5+1) * -1 * atan( 1 / ( -1 + 2^5 ) )   n =  5   d_n = -1-1i 
assign v[4'b1111] [05] = 21'h 1FF7DF;  // -2.0315754229491265 = 2^(6+1) * -1 * atan( 1 / ( -1 + 2^6 ) )   n =  6   d_n = -1-1i 
assign v[4'b1111] [06] = 21'h 1FF7EF;  // -2.0157063741697390 = 2^(7+1) * -1 * atan( 1 / ( -1 + 2^7 ) )   n =  7   d_n = -1-1i 
assign v[4'b1111] [07] = 21'h 1FF7F7;  // -2.0078328446771208 = 2^(8+1) * -1 * atan( 1 / ( -1 + 2^8 ) )   n =  8   d_n = -1-1i 
assign v[4'b1111] [08] = 21'h 1FF7FB;  // -2.0039113362396619 = 2^(9+1) * -1 * atan( 1 / ( -1 + 2^9 ) )   n =  9   d_n = -1-1i 
assign v[4'b1111] [09] = 21'h 1FF7FD;  // -2.0019543965642979 = 2^(10+1) * -1 * atan( 1 / ( -1 + 2^10 ) )   n = 10   d_n = -1-1i 
assign v[4'b1111] [10] = 21'h 1FF7FE;  // -2.0009768803913479 = 2^(11+1) * -1 * atan( 1 / ( -1 + 2^11 ) )   n = 11   d_n = -1-1i 
assign v[4'b1111] [11] = 21'h 1FF7FF;  // -2.0004883607228541 = 2^(12+1) * -1 * atan( 1 / ( -1 + 2^12 ) )   n = 12   d_n = -1-1i 
assign v[4'b1111] [12] = 21'h 1FF7FF;  // -2.0002441604932146 = 2^(13+1) * -1 * atan( 1 / ( -1 + 2^13 ) )   n = 13   d_n = -1-1i 
assign v[4'b1111] [13] = 21'h 1FF7FF;  // -2.0001220752795539 = 2^(14+1) * -1 * atan( 1 / ( -1 + 2^14 ) )   n = 14   d_n = -1-1i 
assign v[4'b1111] [14] = 21'h 1FF7FF;  // -2.0000610363980136 = 2^(15+1) * -1 * atan( 1 / ( -1 + 2^15 ) )   n = 15   d_n = -1-1i 
assign v[4'b1111] [15] = 21'h 1FF7FF;  // -2.0000305178885660 = 2^(16+1) * -1 * atan( 1 / ( -1 + 2^16 ) )   n = 16   d_n = -1-1i 
assign v[4'b1111] [16] = 21'h 1FF7FF;  // -2.0000152588666729 = 2^(17+1) * -1 * atan( 1 / ( -1 + 2^17 ) )   n = 17   d_n = -1-1i 
assign v[4'b1111] [17] = 21'h 1FF7FF;  // -2.0000076294139340 = 2^(18+1) * -1 * atan( 1 / ( -1 + 2^18 ) )   n = 18   d_n = -1-1i 
assign v[4'b1111] [18] = 21'h 1FF7FF;  // -2.0000038147021164 = 2^(19+1) * -1 * atan( 1 / ( -1 + 2^19 ) )   n = 19   d_n = -1-1i 
assign v[4'b1111] [19] = 21'h 1FF7FF;  // -2.0000019073498456 = 2^(20+1) * -1 * atan( 1 / ( -1 + 2^20 ) )   n = 20   d_n = -1-1i 
assign v[4'b1111] [20] = 21'h 1FF7FF;  // -2.0000009536746197 = 2^(21+1) * -1 * atan( 1 / ( -1 + 2^21 ) )   n = 21   d_n = -1-1i 
assign v[4'b1111] [21] = 21'h 1FF7FF;  // -2.0000004768372341 = 2^(22+1) * -1 * atan( 1 / ( -1 + 2^22 ) )   n = 22   d_n = -1-1i 
assign v[4'b1111] [22] = 21'h 1FF7FF;  // -2.0000002384185982 = 2^(23+1) * -1 * atan( 1 / ( -1 + 2^23 ) )   n = 23   d_n = -1-1i 
assign v[4'b1111] [23] = 21'h 1FF7FF;  // -2.0000001192092944 = 2^(24+1) * -1 * atan( 1 / ( -1 + 2^24 ) )   n = 24   d_n = -1-1i 
assign v[4'b1111] [24] = 21'h 1FF7FF;  // -2.0000000596046461 = 2^(25+1) * -1 * atan( 1 / ( -1 + 2^25 ) )   n = 25   d_n = -1-1i 
assign v[4'b1111] [25] = 21'h 1FF7FF;  // -2.0000000298023228 = 2^(26+1) * -1 * atan( 1 / ( -1 + 2^26 ) )   n = 26   d_n = -1-1i 
assign v[4'b1111] [26] = 21'h 1FF7FF;  // -2.0000000149011612 = 2^(27+1) * -1 * atan( 1 / ( -1 + 2^27 ) )   n = 27   d_n = -1-1i 
assign v[4'b1111] [27] = 21'h 1FF7FF;  // -2.0000000074505806 = 2^(28+1) * -1 * atan( 1 / ( -1 + 2^28 ) )   n = 28   d_n = -1-1i 
assign v[4'b1111] [28] = 21'h 1FF7FF;  // -2.0000000037252903 = 2^(29+1) * -1 * atan( 1 / ( -1 + 2^29 ) )   n = 29   d_n = -1-1i 
assign v[4'b1111] [29] = 21'h 1FF7FF;  // -2.0000000018626451 = 2^(30+1) * -1 * atan( 1 / ( -1 + 2^30 ) )   n = 30   d_n = -1-1i 
assign v[4'b1111] [30] = 21'h 1FF7FF;  // -2.0000000009313226 = 2^(31+1) * -1 * atan( 1 / ( -1 + 2^31 ) )   n = 31   d_n = -1-1i 
assign v[4'b1111] [31] = 21'h 1FF7FF;  // -2.0000000004656613 = 2^(32+1) * -1 * atan( 1 / ( -1 + 2^32 ) )   n = 32   d_n = -1-1i 
assign v[4'b1111] [32] = 21'h 1FF7FF;  // -2.0000000002328306 = 2^(33+1) * -1 * atan( 1 / ( -1 + 2^33 ) )   n = 33   d_n = -1-1i 
assign v[4'b1111] [33] = 21'h 1FF7FF;  // -2.0000000001164153 = 2^(34+1) * -1 * atan( 1 / ( -1 + 2^34 ) )   n = 34   d_n = -1-1i 
assign v[4'b1111] [34] = 21'h 1FF7FF;  // -2.0000000000582077 = 2^(35+1) * -1 * atan( 1 / ( -1 + 2^35 ) )   n = 35   d_n = -1-1i 
assign v[4'b1111] [35] = 21'h 1FF7FF;  // -2.0000000000291038 = 2^(36+1) * -1 * atan( 1 / ( -1 + 2^36 ) )   n = 36   d_n = -1-1i 
assign v[4'b1111] [36] = 21'h 1FF7FF;  // -2.0000000000145519 = 2^(37+1) * -1 * atan( 1 / ( -1 + 2^37 ) )   n = 37   d_n = -1-1i 
assign v[4'b1111] [37] = 21'h 1FF7FF;  // -2.0000000000072760 = 2^(38+1) * -1 * atan( 1 / ( -1 + 2^38 ) )   n = 38   d_n = -1-1i 
assign v[4'b1111] [38] = 21'h 1FF7FF;  // -2.0000000000036380 = 2^(39+1) * -1 * atan( 1 / ( -1 + 2^39 ) )   n = 39   d_n = -1-1i 
assign v[4'b1111] [39] = 21'h 1FF7FF;  // -2.0000000000018190 = 2^(40+1) * -1 * atan( 1 / ( -1 + 2^40 ) )   n = 40   d_n = -1-1i 
assign v[4'b1111] [40] = 21'h 1FF7FF;  // -2.0000000000009095 = 2^(41+1) * -1 * atan( 1 / ( -1 + 2^41 ) )   n = 41   d_n = -1-1i 
assign v[4'b1111] [41] = 21'h 1FF7FF;  // -2.0000000000004547 = 2^(42+1) * -1 * atan( 1 / ( -1 + 2^42 ) )   n = 42   d_n = -1-1i 
assign v[4'b1111] [42] = 21'h 1FF7FF;  // -2.0000000000002274 = 2^(43+1) * -1 * atan( 1 / ( -1 + 2^43 ) )   n = 43   d_n = -1-1i 
assign v[4'b1111] [43] = 21'h 1FF800;  // -2.0000000000001137 = 2^(44+1) * -1 * atan( 1 / ( -1 + 2^44 ) )   n = 44   d_n = -1-1i 
assign v[4'b1111] [44] = 21'h 1FF800;  // -2.0000000000000568 = 2^(45+1) * -1 * atan( 1 / ( -1 + 2^45 ) )   n = 45   d_n = -1-1i 
assign v[4'b1111] [45] = 21'h 1FF800;  // -2.0000000000000284 = 2^(46+1) * -1 * atan( 1 / ( -1 + 2^46 ) )   n = 46   d_n = -1-1i 
assign v[4'b1111] [46] = 21'h 1FF800;  // -2.0000000000000142 = 2^(47+1) * -1 * atan( 1 / ( -1 + 2^47 ) )   n = 47   d_n = -1-1i 
assign v[4'b1111] [47] = 21'h 1FF800;  // -2.0000000000000071 = 2^(48+1) * -1 * atan( 1 / ( -1 + 2^48 ) )   n = 48   d_n = -1-1i 
assign v[4'b1111] [48] = 21'h 1FF800;  // -2.0000000000000036 = 2^(49+1) * -1 * atan( 1 / ( -1 + 2^49 ) )   n = 49   d_n = -1-1i 
assign v[4'b1111] [49] = 21'h 1FF800;  // -2.0000000000000018 = 2^(50+1) * -1 * atan( 1 / ( -1 + 2^50 ) )   n = 50   d_n = -1-1i 
assign v[4'b1111] [50] = 21'h 1FF800;  // -2.0000000000000009 = 2^(51+1) * -1 * atan( 1 / ( -1 + 2^51 ) )   n = 51   d_n = -1-1i 
assign v[4'b1111] [51] = 21'h 1FF800;  // -2.0000000000000004 = 2^(52+1) * -1 * atan( 1 / ( -1 + 2^52 ) )   n = 52   d_n = -1-1i 
assign v[4'b1111] [52] = 21'h 1FF800;  // -2.0000000000000004 = 2^(53+1) * -1 * atan( 1 / ( -1 + 2^53 ) )   n = 53   d_n = -1-1i 
assign v[4'b1111] [53] = 21'h 1FF800;  // -2.0000000000000000 = 2^(54+1) * -1 * atan( 1 / ( -1 + 2^54 ) )   n = 54   d_n = -1-1i 
assign v[4'b1111] [54] = 21'h 1FF800;  // -2.0000000000000000 = 2^(55+1) * -1 * atan( 1 / ( -1 + 2^55 ) )   n = 55   d_n = -1-1i 
assign v[4'b1111] [55] = 21'h 1FF800;  // -2.0000000000000000 = 2^(56+1) * -1 * atan( 1 / ( -1 + 2^56 ) )   n = 56   d_n = -1-1i 
assign v[4'b1111] [56] = 21'h 1FF800;  // -2.0000000000000000 = 2^(57+1) * -1 * atan( 1 / ( -1 + 2^57 ) )   n = 57   d_n = -1-1i 
assign v[4'b1111] [57] = 21'h 1FF800;  // -2.0000000000000000 = 2^(58+1) * -1 * atan( 1 / ( -1 + 2^58 ) )   n = 58   d_n = -1-1i 
assign v[4'b1111] [58] = 21'h 1FF800;  // -2.0000000000000000 = 2^(59+1) * -1 * atan( 1 / ( -1 + 2^59 ) )   n = 59   d_n = -1-1i 
assign v[4'b1111] [59] = 21'h 1FF800;  // -2.0000000000000000 = 2^(60+1) * -1 * atan( 1 / ( -1 + 2^60 ) )   n = 60   d_n = -1-1i 
assign v[4'b1111] [60] = 21'h 1FF800;  // -2.0000000000000000 = 2^(61+1) * -1 * atan( 1 / ( -1 + 2^61 ) )   n = 61   d_n = -1-1i 
assign v[4'b1111] [61] = 21'h 1FF800;  // -2.0000000000000000 = 2^(62+1) * -1 * atan( 1 / ( -1 + 2^62 ) )   n = 62   d_n = -1-1i 
assign v[4'b1111] [62] = 21'h 1FF800;  // -2.0000000000000000 = 2^(63+1) * -1 * atan( 1 / ( -1 + 2^63 ) )   n = 63   d_n = -1-1i 
assign v[4'b1111] [63] = 21'h 1FF800;  // -2.0000000000000000 = 2^(64+1) * -1 * atan( 1 / ( -1 + 2^64 ) )   n = 64   d_n = -1-1i 
