// -----------------------------------------------------------------------------
//  Copyright (c) 2016 Microelectronics Lab. FIUBA.
//  All Rights Reserved.
//
//  The information contained in this file is confidential and proprietary.
//  Any reproduction, use or disclosure, in whole or in part, of this
//  program, including any attempt to obtain a human-readable version of this
//  program, without the express, prior written consent of Microelectronics Lab.
//  FIUBA is strictly prohibited.
//
// -----------------------------------------------------------------------------
// Description:
// ------------
//
// Monitor for lut_decoder block.
//
// -----------------------------------------------------------------------------
// File name:
// ----------
//
// lut_decoder_monitor.v
//
// -----------------------------------------------------------------------------
// History:
// --------
//
//    - 2016-08-28 - ilesser - Initial version.
//
// -----------------------------------------------------------------------------

`include "/home/ilesser/simlib/simlib_defs.vh"

// *****************************************************************************
// Interface
// *****************************************************************************
module lut_decoder_monitor #(
   // ----------------------------------
   // Parameters
   // ----------------------------------
   parameter W       = 64
   ) (
   // ----------------------------------
   // Clock, reset & enable inputs
   // ----------------------------------
   input wire              clk,
   input wire              arst,
   input wire              srst,
   input wire              enable,
   // ----------------------------------
   // Data inputs
   // ----------------------------------
   input  wire [2*W-1:0]   lut_X_n_csd,
   input  wire [2*W-1:0]   lut_Y_n_csd,
   // ----------------------------------
   // Data outputs
   // ----------------------------------
   output wire [W-1:0]     res_lut_X_n,
   output wire [W-1:0]     res_lut_Y_n
   );
// *****************************************************************************

// *****************************************************************************
// Architecture
// *****************************************************************************

   // -----------------------------------------------------
   // Internal signals
   // -----------------------------------------------------
   // -----------------------------------------------------

   csd2bin #(
    // ----------------------------------
    // Parameters
    // ----------------------------------
      .W                   (W)
   ) csd2bin_X (
    // ----------------------------------
    // Data inputs
    // ----------------------------------
      .x                   (lut_X_n_csd),
    // ----------------------------------
    // Data outputs
    // ----------------------------------
      .y                   (res_lut_X_n)
   );

   csd2bin #(
    // ----------------------------------
    // Parameters
    // ----------------------------------
      .W                   (W)
   ) csd2bin_Y (
    // ----------------------------------
    // Data inputs
    // ----------------------------------
      .x                   (lut_Y_n_csd),
    // ----------------------------------
    // Data outputs
    // ----------------------------------
      .y                   (res_lut_Y_n)
   );
// *****************************************************************************

`ifdef RTL_DEBUG

//

`else

//XXXXX FILL IN HERE XXXXX

`endif
// *****************************************************************************

endmodule



