assign X[4'b0000] [01] = 64'h0000000000000000;
assign Y[4'b0000] [01] = 64'h00000000000003C0;
assign u[4'b0000] [01] = 64'h00000000000007C0;
assign v[4'b0000] [01] = 64'h0000000000000BC0;
assign X[4'b0000] [02] = 64'h0000000000000001;
assign Y[4'b0000] [02] = 64'h00000000000003C1;
assign u[4'b0000] [02] = 64'h00000000000007C1;
assign v[4'b0000] [02] = 64'h0000000000000BC1;
assign X[4'b0000] [03] = 64'h0000000000000002;
assign Y[4'b0000] [03] = 64'h00000000000003C2;
assign u[4'b0000] [03] = 64'h00000000000007C2;
assign v[4'b0000] [03] = 64'h0000000000000BC2;
assign X[4'b0000] [04] = 64'h0000000000000003;
assign Y[4'b0000] [04] = 64'h00000000000003C3;
assign u[4'b0000] [04] = 64'h00000000000007C3;
assign v[4'b0000] [04] = 64'h0000000000000BC3;
assign X[4'b0000] [05] = 64'h0000000000000004;
assign Y[4'b0000] [05] = 64'h00000000000003C4;
assign u[4'b0000] [05] = 64'h00000000000007C4;
assign v[4'b0000] [05] = 64'h0000000000000BC4;
assign X[4'b0000] [06] = 64'h0000000000000005;
assign Y[4'b0000] [06] = 64'h00000000000003C5;
assign u[4'b0000] [06] = 64'h00000000000007C5;
assign v[4'b0000] [06] = 64'h0000000000000BC5;
assign X[4'b0000] [07] = 64'h0000000000000006;
assign Y[4'b0000] [07] = 64'h00000000000003C6;
assign u[4'b0000] [07] = 64'h00000000000007C6;
assign v[4'b0000] [07] = 64'h0000000000000BC6;
assign X[4'b0000] [08] = 64'h0000000000000007;
assign Y[4'b0000] [08] = 64'h00000000000003C7;
assign u[4'b0000] [08] = 64'h00000000000007C7;
assign v[4'b0000] [08] = 64'h0000000000000BC7;
assign X[4'b0000] [09] = 64'h0000000000000008;
assign Y[4'b0000] [09] = 64'h00000000000003C8;
assign u[4'b0000] [09] = 64'h00000000000007C8;
assign v[4'b0000] [09] = 64'h0000000000000BC8;
assign X[4'b0000] [10] = 64'h0000000000000009;
assign Y[4'b0000] [10] = 64'h00000000000003C9;
assign u[4'b0000] [10] = 64'h00000000000007C9;
assign v[4'b0000] [10] = 64'h0000000000000BC9;
assign X[4'b0000] [11] = 64'h000000000000000A;
assign Y[4'b0000] [11] = 64'h00000000000003CA;
assign u[4'b0000] [11] = 64'h00000000000007CA;
assign v[4'b0000] [11] = 64'h0000000000000BCA;
assign X[4'b0000] [12] = 64'h000000000000000B;
assign Y[4'b0000] [12] = 64'h00000000000003CB;
assign u[4'b0000] [12] = 64'h00000000000007CB;
assign v[4'b0000] [12] = 64'h0000000000000BCB;
assign X[4'b0000] [13] = 64'h000000000000000C;
assign Y[4'b0000] [13] = 64'h00000000000003CC;
assign u[4'b0000] [13] = 64'h00000000000007CC;
assign v[4'b0000] [13] = 64'h0000000000000BCC;
assign X[4'b0000] [14] = 64'h000000000000000D;
assign Y[4'b0000] [14] = 64'h00000000000003CD;
assign u[4'b0000] [14] = 64'h00000000000007CD;
assign v[4'b0000] [14] = 64'h0000000000000BCD;
assign X[4'b0000] [15] = 64'h000000000000000E;
assign Y[4'b0000] [15] = 64'h00000000000003CE;
assign u[4'b0000] [15] = 64'h00000000000007CE;
assign v[4'b0000] [15] = 64'h0000000000000BCE;
assign X[4'b0000] [16] = 64'h000000000000000F;
assign Y[4'b0000] [16] = 64'h00000000000003CF;
assign u[4'b0000] [16] = 64'h00000000000007CF;
assign v[4'b0000] [16] = 64'h0000000000000BCF;
assign X[4'b0000] [17] = 64'h0000000000000010;
assign Y[4'b0000] [17] = 64'h00000000000003D0;
assign u[4'b0000] [17] = 64'h00000000000007D0;
assign v[4'b0000] [17] = 64'h0000000000000BD0;
assign X[4'b0000] [18] = 64'h0000000000000011;
assign Y[4'b0000] [18] = 64'h00000000000003D1;
assign u[4'b0000] [18] = 64'h00000000000007D1;
assign v[4'b0000] [18] = 64'h0000000000000BD1;
assign X[4'b0000] [19] = 64'h0000000000000012;
assign Y[4'b0000] [19] = 64'h00000000000003D2;
assign u[4'b0000] [19] = 64'h00000000000007D2;
assign v[4'b0000] [19] = 64'h0000000000000BD2;
assign X[4'b0000] [20] = 64'h0000000000000013;
assign Y[4'b0000] [20] = 64'h00000000000003D3;
assign u[4'b0000] [20] = 64'h00000000000007D3;
assign v[4'b0000] [20] = 64'h0000000000000BD3;
assign X[4'b0000] [21] = 64'h0000000000000014;
assign Y[4'b0000] [21] = 64'h00000000000003D4;
assign u[4'b0000] [21] = 64'h00000000000007D4;
assign v[4'b0000] [21] = 64'h0000000000000BD4;
assign X[4'b0000] [22] = 64'h0000000000000015;
assign Y[4'b0000] [22] = 64'h00000000000003D5;
assign u[4'b0000] [22] = 64'h00000000000007D5;
assign v[4'b0000] [22] = 64'h0000000000000BD5;
assign X[4'b0000] [23] = 64'h0000000000000016;
assign Y[4'b0000] [23] = 64'h00000000000003D6;
assign u[4'b0000] [23] = 64'h00000000000007D6;
assign v[4'b0000] [23] = 64'h0000000000000BD6;
assign X[4'b0000] [24] = 64'h0000000000000017;
assign Y[4'b0000] [24] = 64'h00000000000003D7;
assign u[4'b0000] [24] = 64'h00000000000007D7;
assign v[4'b0000] [24] = 64'h0000000000000BD7;
assign X[4'b0000] [25] = 64'h0000000000000018;
assign Y[4'b0000] [25] = 64'h00000000000003D8;
assign u[4'b0000] [25] = 64'h00000000000007D8;
assign v[4'b0000] [25] = 64'h0000000000000BD8;
assign X[4'b0000] [26] = 64'h0000000000000019;
assign Y[4'b0000] [26] = 64'h00000000000003D9;
assign u[4'b0000] [26] = 64'h00000000000007D9;
assign v[4'b0000] [26] = 64'h0000000000000BD9;
assign X[4'b0000] [27] = 64'h000000000000001A;
assign Y[4'b0000] [27] = 64'h00000000000003DA;
assign u[4'b0000] [27] = 64'h00000000000007DA;
assign v[4'b0000] [27] = 64'h0000000000000BDA;
assign X[4'b0000] [28] = 64'h000000000000001B;
assign Y[4'b0000] [28] = 64'h00000000000003DB;
assign u[4'b0000] [28] = 64'h00000000000007DB;
assign v[4'b0000] [28] = 64'h0000000000000BDB;
assign X[4'b0000] [29] = 64'h000000000000001C;
assign Y[4'b0000] [29] = 64'h00000000000003DC;
assign u[4'b0000] [29] = 64'h00000000000007DC;
assign v[4'b0000] [29] = 64'h0000000000000BDC;
assign X[4'b0000] [30] = 64'h000000000000001D;
assign Y[4'b0000] [30] = 64'h00000000000003DD;
assign u[4'b0000] [30] = 64'h00000000000007DD;
assign v[4'b0000] [30] = 64'h0000000000000BDD;
assign X[4'b0000] [31] = 64'h000000000000001E;
assign Y[4'b0000] [31] = 64'h00000000000003DE;
assign u[4'b0000] [31] = 64'h00000000000007DE;
assign v[4'b0000] [31] = 64'h0000000000000BDE;
assign X[4'b0000] [32] = 64'h000000000000001F;
assign Y[4'b0000] [32] = 64'h00000000000003DF;
assign u[4'b0000] [32] = 64'h00000000000007DF;
assign v[4'b0000] [32] = 64'h0000000000000BDF;
assign X[4'b0000] [33] = 64'h0000000000000020;
assign Y[4'b0000] [33] = 64'h00000000000003E0;
assign u[4'b0000] [33] = 64'h00000000000007E0;
assign v[4'b0000] [33] = 64'h0000000000000BE0;
assign X[4'b0000] [34] = 64'h0000000000000021;
assign Y[4'b0000] [34] = 64'h00000000000003E1;
assign u[4'b0000] [34] = 64'h00000000000007E1;
assign v[4'b0000] [34] = 64'h0000000000000BE1;
assign X[4'b0000] [35] = 64'h0000000000000022;
assign Y[4'b0000] [35] = 64'h00000000000003E2;
assign u[4'b0000] [35] = 64'h00000000000007E2;
assign v[4'b0000] [35] = 64'h0000000000000BE2;
assign X[4'b0000] [36] = 64'h0000000000000023;
assign Y[4'b0000] [36] = 64'h00000000000003E3;
assign u[4'b0000] [36] = 64'h00000000000007E3;
assign v[4'b0000] [36] = 64'h0000000000000BE3;
assign X[4'b0000] [37] = 64'h0000000000000024;
assign Y[4'b0000] [37] = 64'h00000000000003E4;
assign u[4'b0000] [37] = 64'h00000000000007E4;
assign v[4'b0000] [37] = 64'h0000000000000BE4;
assign X[4'b0000] [38] = 64'h0000000000000025;
assign Y[4'b0000] [38] = 64'h00000000000003E5;
assign u[4'b0000] [38] = 64'h00000000000007E5;
assign v[4'b0000] [38] = 64'h0000000000000BE5;
assign X[4'b0000] [39] = 64'h0000000000000026;
assign Y[4'b0000] [39] = 64'h00000000000003E6;
assign u[4'b0000] [39] = 64'h00000000000007E6;
assign v[4'b0000] [39] = 64'h0000000000000BE6;
assign X[4'b0000] [40] = 64'h0000000000000027;
assign Y[4'b0000] [40] = 64'h00000000000003E7;
assign u[4'b0000] [40] = 64'h00000000000007E7;
assign v[4'b0000] [40] = 64'h0000000000000BE7;
assign X[4'b0000] [41] = 64'h0000000000000028;
assign Y[4'b0000] [41] = 64'h00000000000003E8;
assign u[4'b0000] [41] = 64'h00000000000007E8;
assign v[4'b0000] [41] = 64'h0000000000000BE8;
assign X[4'b0000] [42] = 64'h0000000000000029;
assign Y[4'b0000] [42] = 64'h00000000000003E9;
assign u[4'b0000] [42] = 64'h00000000000007E9;
assign v[4'b0000] [42] = 64'h0000000000000BE9;
assign X[4'b0000] [43] = 64'h000000000000002A;
assign Y[4'b0000] [43] = 64'h00000000000003EA;
assign u[4'b0000] [43] = 64'h00000000000007EA;
assign v[4'b0000] [43] = 64'h0000000000000BEA;
assign X[4'b0000] [44] = 64'h000000000000002B;
assign Y[4'b0000] [44] = 64'h00000000000003EB;
assign u[4'b0000] [44] = 64'h00000000000007EB;
assign v[4'b0000] [44] = 64'h0000000000000BEB;
assign X[4'b0000] [45] = 64'h000000000000002C;
assign Y[4'b0000] [45] = 64'h00000000000003EC;
assign u[4'b0000] [45] = 64'h00000000000007EC;
assign v[4'b0000] [45] = 64'h0000000000000BEC;
assign X[4'b0000] [46] = 64'h000000000000002D;
assign Y[4'b0000] [46] = 64'h00000000000003ED;
assign u[4'b0000] [46] = 64'h00000000000007ED;
assign v[4'b0000] [46] = 64'h0000000000000BED;
assign X[4'b0000] [47] = 64'h000000000000002E;
assign Y[4'b0000] [47] = 64'h00000000000003EE;
assign u[4'b0000] [47] = 64'h00000000000007EE;
assign v[4'b0000] [47] = 64'h0000000000000BEE;
assign X[4'b0000] [48] = 64'h000000000000002F;
assign Y[4'b0000] [48] = 64'h00000000000003EF;
assign u[4'b0000] [48] = 64'h00000000000007EF;
assign v[4'b0000] [48] = 64'h0000000000000BEF;
assign X[4'b0000] [49] = 64'h0000000000000030;
assign Y[4'b0000] [49] = 64'h00000000000003F0;
assign u[4'b0000] [49] = 64'h00000000000007F0;
assign v[4'b0000] [49] = 64'h0000000000000BF0;
assign X[4'b0000] [50] = 64'h0000000000000031;
assign Y[4'b0000] [50] = 64'h00000000000003F1;
assign u[4'b0000] [50] = 64'h00000000000007F1;
assign v[4'b0000] [50] = 64'h0000000000000BF1;
assign X[4'b0000] [51] = 64'h0000000000000032;
assign Y[4'b0000] [51] = 64'h00000000000003F2;
assign u[4'b0000] [51] = 64'h00000000000007F2;
assign v[4'b0000] [51] = 64'h0000000000000BF2;
assign X[4'b0000] [52] = 64'h0000000000000033;
assign Y[4'b0000] [52] = 64'h00000000000003F3;
assign u[4'b0000] [52] = 64'h00000000000007F3;
assign v[4'b0000] [52] = 64'h0000000000000BF3;
assign X[4'b0000] [53] = 64'h0000000000000034;
assign Y[4'b0000] [53] = 64'h00000000000003F4;
assign u[4'b0000] [53] = 64'h00000000000007F4;
assign v[4'b0000] [53] = 64'h0000000000000BF4;
assign X[4'b0000] [54] = 64'h0000000000000035;
assign Y[4'b0000] [54] = 64'h00000000000003F5;
assign u[4'b0000] [54] = 64'h00000000000007F5;
assign v[4'b0000] [54] = 64'h0000000000000BF5;
assign X[4'b0000] [55] = 64'h0000000000000036;
assign Y[4'b0000] [55] = 64'h00000000000003F6;
assign u[4'b0000] [55] = 64'h00000000000007F6;
assign v[4'b0000] [55] = 64'h0000000000000BF6;
assign X[4'b0000] [56] = 64'h0000000000000037;
assign Y[4'b0000] [56] = 64'h00000000000003F7;
assign u[4'b0000] [56] = 64'h00000000000007F7;
assign v[4'b0000] [56] = 64'h0000000000000BF7;
assign X[4'b0000] [57] = 64'h0000000000000038;
assign Y[4'b0000] [57] = 64'h00000000000003F8;
assign u[4'b0000] [57] = 64'h00000000000007F8;
assign v[4'b0000] [57] = 64'h0000000000000BF8;
assign X[4'b0000] [58] = 64'h0000000000000039;
assign Y[4'b0000] [58] = 64'h00000000000003F9;
assign u[4'b0000] [58] = 64'h00000000000007F9;
assign v[4'b0000] [58] = 64'h0000000000000BF9;
assign X[4'b0000] [59] = 64'h000000000000003A;
assign Y[4'b0000] [59] = 64'h00000000000003FA;
assign u[4'b0000] [59] = 64'h00000000000007FA;
assign v[4'b0000] [59] = 64'h0000000000000BFA;
assign X[4'b0000] [60] = 64'h000000000000003B;
assign Y[4'b0000] [60] = 64'h00000000000003FB;
assign u[4'b0000] [60] = 64'h00000000000007FB;
assign v[4'b0000] [60] = 64'h0000000000000BFB;
assign X[4'b0000] [61] = 64'h000000000000003C;
assign Y[4'b0000] [61] = 64'h00000000000003FC;
assign u[4'b0000] [61] = 64'h00000000000007FC;
assign v[4'b0000] [61] = 64'h0000000000000BFC;
assign X[4'b0000] [62] = 64'h000000000000003D;
assign Y[4'b0000] [62] = 64'h00000000000003FD;
assign u[4'b0000] [62] = 64'h00000000000007FD;
assign v[4'b0000] [62] = 64'h0000000000000BFD;
assign X[4'b0000] [63] = 64'h000000000000003E;
assign Y[4'b0000] [63] = 64'h00000000000003FE;
assign u[4'b0000] [63] = 64'h00000000000007FE;
assign v[4'b0000] [63] = 64'h0000000000000BFE;
assign X[4'b0000] [64] = 64'h000000000000003F;
assign Y[4'b0000] [64] = 64'h00000000000003FF;
assign u[4'b0000] [64] = 64'h00000000000007FF;
assign v[4'b0000] [64] = 64'h0000000000000BFF;
assign X[4'b0001] [01] = 64'h0000000000000040;
assign Y[4'b0001] [01] = 64'h0000000000000400;
assign u[4'b0001] [01] = 64'h0000000000000800;
assign v[4'b0001] [01] = 64'h0000000000000C00;
assign X[4'b0001] [02] = 64'h0000000000000041;
assign Y[4'b0001] [02] = 64'h0000000000000401;
assign u[4'b0001] [02] = 64'h0000000000000801;
assign v[4'b0001] [02] = 64'h0000000000000C01;
assign X[4'b0001] [03] = 64'h0000000000000042;
assign Y[4'b0001] [03] = 64'h0000000000000402;
assign u[4'b0001] [03] = 64'h0000000000000802;
assign v[4'b0001] [03] = 64'h0000000000000C02;
assign X[4'b0001] [04] = 64'h0000000000000043;
assign Y[4'b0001] [04] = 64'h0000000000000403;
assign u[4'b0001] [04] = 64'h0000000000000803;
assign v[4'b0001] [04] = 64'h0000000000000C03;
assign X[4'b0001] [05] = 64'h0000000000000044;
assign Y[4'b0001] [05] = 64'h0000000000000404;
assign u[4'b0001] [05] = 64'h0000000000000804;
assign v[4'b0001] [05] = 64'h0000000000000C04;
assign X[4'b0001] [06] = 64'h0000000000000045;
assign Y[4'b0001] [06] = 64'h0000000000000405;
assign u[4'b0001] [06] = 64'h0000000000000805;
assign v[4'b0001] [06] = 64'h0000000000000C05;
assign X[4'b0001] [07] = 64'h0000000000000046;
assign Y[4'b0001] [07] = 64'h0000000000000406;
assign u[4'b0001] [07] = 64'h0000000000000806;
assign v[4'b0001] [07] = 64'h0000000000000C06;
assign X[4'b0001] [08] = 64'h0000000000000047;
assign Y[4'b0001] [08] = 64'h0000000000000407;
assign u[4'b0001] [08] = 64'h0000000000000807;
assign v[4'b0001] [08] = 64'h0000000000000C07;
assign X[4'b0001] [09] = 64'h0000000000000048;
assign Y[4'b0001] [09] = 64'h0000000000000408;
assign u[4'b0001] [09] = 64'h0000000000000808;
assign v[4'b0001] [09] = 64'h0000000000000C08;
assign X[4'b0001] [10] = 64'h0000000000000049;
assign Y[4'b0001] [10] = 64'h0000000000000409;
assign u[4'b0001] [10] = 64'h0000000000000809;
assign v[4'b0001] [10] = 64'h0000000000000C09;
assign X[4'b0001] [11] = 64'h000000000000004A;
assign Y[4'b0001] [11] = 64'h000000000000040A;
assign u[4'b0001] [11] = 64'h000000000000080A;
assign v[4'b0001] [11] = 64'h0000000000000C0A;
assign X[4'b0001] [12] = 64'h000000000000004B;
assign Y[4'b0001] [12] = 64'h000000000000040B;
assign u[4'b0001] [12] = 64'h000000000000080B;
assign v[4'b0001] [12] = 64'h0000000000000C0B;
assign X[4'b0001] [13] = 64'h000000000000004C;
assign Y[4'b0001] [13] = 64'h000000000000040C;
assign u[4'b0001] [13] = 64'h000000000000080C;
assign v[4'b0001] [13] = 64'h0000000000000C0C;
assign X[4'b0001] [14] = 64'h000000000000004D;
assign Y[4'b0001] [14] = 64'h000000000000040D;
assign u[4'b0001] [14] = 64'h000000000000080D;
assign v[4'b0001] [14] = 64'h0000000000000C0D;
assign X[4'b0001] [15] = 64'h000000000000004E;
assign Y[4'b0001] [15] = 64'h000000000000040E;
assign u[4'b0001] [15] = 64'h000000000000080E;
assign v[4'b0001] [15] = 64'h0000000000000C0E;
assign X[4'b0001] [16] = 64'h000000000000004F;
assign Y[4'b0001] [16] = 64'h000000000000040F;
assign u[4'b0001] [16] = 64'h000000000000080F;
assign v[4'b0001] [16] = 64'h0000000000000C0F;
assign X[4'b0001] [17] = 64'h0000000000000050;
assign Y[4'b0001] [17] = 64'h0000000000000410;
assign u[4'b0001] [17] = 64'h0000000000000810;
assign v[4'b0001] [17] = 64'h0000000000000C10;
assign X[4'b0001] [18] = 64'h0000000000000051;
assign Y[4'b0001] [18] = 64'h0000000000000411;
assign u[4'b0001] [18] = 64'h0000000000000811;
assign v[4'b0001] [18] = 64'h0000000000000C11;
assign X[4'b0001] [19] = 64'h0000000000000052;
assign Y[4'b0001] [19] = 64'h0000000000000412;
assign u[4'b0001] [19] = 64'h0000000000000812;
assign v[4'b0001] [19] = 64'h0000000000000C12;
assign X[4'b0001] [20] = 64'h0000000000000053;
assign Y[4'b0001] [20] = 64'h0000000000000413;
assign u[4'b0001] [20] = 64'h0000000000000813;
assign v[4'b0001] [20] = 64'h0000000000000C13;
assign X[4'b0001] [21] = 64'h0000000000000054;
assign Y[4'b0001] [21] = 64'h0000000000000414;
assign u[4'b0001] [21] = 64'h0000000000000814;
assign v[4'b0001] [21] = 64'h0000000000000C14;
assign X[4'b0001] [22] = 64'h0000000000000055;
assign Y[4'b0001] [22] = 64'h0000000000000415;
assign u[4'b0001] [22] = 64'h0000000000000815;
assign v[4'b0001] [22] = 64'h0000000000000C15;
assign X[4'b0001] [23] = 64'h0000000000000056;
assign Y[4'b0001] [23] = 64'h0000000000000416;
assign u[4'b0001] [23] = 64'h0000000000000816;
assign v[4'b0001] [23] = 64'h0000000000000C16;
assign X[4'b0001] [24] = 64'h0000000000000000;
assign X[4'b0010] [47] = 64'h00000000000000AE;
assign X[4'b0010] [48] = 64'h0000000000000000;
assign X[4'b0010] [48] = 64'h00000000000000AF;
assign X[4'b0010] [49] = 64'h0000000000000000;
assign X[4'b0010] [49] = 64'h00000000000000B0;
assign X[4'b0010] [50] = 64'h0000000000000000;
assign X[4'b0010] [50] = 64'h00000000000000B1;
assign X[4'b0010] [51] = 64'h0000000000000000;
assign X[4'b0010] [51] = 64'h00000000000000B2;
assign X[4'b0010] [52] = 64'h0000000000000000;
assign X[4'b0010] [52] = 64'h00000000000000B3;
assign X[4'b0010] [53] = 64'h0000000000000000;
assign X[4'b0010] [53] = 64'h00000000000000B4;
assign X[4'b0010] [54] = 64'h0000000000000000;
assign X[4'b0010] [54] = 64'h00000000000000B5;
assign X[4'b0010] [55] = 64'h0000000000000000;
assign X[4'b0010] [55] = 64'h00000000000000B6;
assign X[4'b0010] [56] = 64'h0000000000000000;
assign X[4'b0010] [56] = 64'h00000000000000B7;
assign X[4'b0010] [57] = 64'h0000000000000000;
assign X[4'b0010] [57] = 64'h00000000000000B8;
assign X[4'b0010] [58] = 64'h0000000000000000;
assign X[4'b0010] [58] = 64'h00000000000000B9;
assign X[4'b0010] [59] = 64'h0000000000000000;
assign X[4'b0010] [59] = 64'h00000000000000BA;
assign X[4'b0010] [60] = 64'h0000000000000000;
assign X[4'b0010] [60] = 64'h00000000000000BB;
assign X[4'b0010] [61] = 64'h0000000000000000;
assign X[4'b0010] [61] = 64'h00000000000000BC;
assign X[4'b0010] [62] = 64'h0000000000000000;
assign X[4'b0010] [62] = 64'h00000000000000BD;
assign X[4'b0010] [63] = 64'h0000000000000000;
assign X[4'b0010] [63] = 64'h00000000000000BE;
assign X[4'b0010] [64] = 64'h0000000000000000;
assign X[4'b0010] [64] = 64'h00000000000000BF;
assign X[4'b0001] [33] = 64'h0000000000000060;
assign Y[4'b0001] [33] = 64'h0000000000000420;
assign u[4'b0001] [33] = 64'h0000000000000820;
assign v[4'b0001] [33] = 64'h0000000000000C20;
assign X[4'b0001] [34] = 64'h0000000000000061;
assign Y[4'b0001] [34] = 64'h0000000000000421;
assign u[4'b0001] [34] = 64'h0000000000000821;
assign v[4'b0001] [34] = 64'h0000000000000C21;
assign X[4'b0001] [35] = 64'h0000000000000062;
assign Y[4'b0001] [35] = 64'h0000000000000422;
assign u[4'b0001] [35] = 64'h0000000000000822;
assign v[4'b0001] [35] = 64'h0000000000000C22;
assign X[4'b0001] [36] = 64'h0000000000000063;
assign Y[4'b0001] [36] = 64'h0000000000000423;
assign u[4'b0001] [36] = 64'h0000000000000823;
assign v[4'b0001] [36] = 64'h0000000000000C23;
assign X[4'b0001] [37] = 64'h0000000000000064;
assign Y[4'b0001] [37] = 64'h0000000000000424;
assign u[4'b0001] [37] = 64'h0000000000000824;
assign v[4'b0001] [37] = 64'h0000000000000C24;
assign X[4'b0001] [38] = 64'h0000000000000065;
assign Y[4'b0001] [38] = 64'h0000000000000425;
assign u[4'b0001] [38] = 64'h0000000000000825;
assign v[4'b0001] [38] = 64'h0000000000000C25;
assign X[4'b0001] [39] = 64'h0000000000000066;
assign Y[4'b0001] [39] = 64'h0000000000000426;
assign u[4'b0001] [39] = 64'h0000000000000826;
assign v[4'b0001] [39] = 64'h0000000000000C26;
assign X[4'b0001] [40] = 64'h0000000000000067;
assign Y[4'b0001] [40] = 64'h0000000000000427;
assign u[4'b0001] [40] = 64'h0000000000000827;
assign v[4'b0001] [40] = 64'h0000000000000C27;
assign X[4'b0001] [41] = 64'h0000000000000068;
assign Y[4'b0001] [41] = 64'h0000000000000428;
assign u[4'b0001] [41] = 64'h0000000000000828;
assign v[4'b0001] [41] = 64'h0000000000000C28;
assign X[4'b0001] [42] = 64'h0000000000000069;
assign Y[4'b0001] [42] = 64'h0000000000000429;
assign u[4'b0001] [42] = 64'h0000000000000829;
assign v[4'b0001] [42] = 64'h0000000000000C29;
assign X[4'b0001] [43] = 64'h000000000000006A;
assign Y[4'b0001] [43] = 64'h000000000000042A;
assign u[4'b0001] [43] = 64'h000000000000082A;
assign v[4'b0001] [43] = 64'h0000000000000C2A;
assign X[4'b0001] [44] = 64'h000000000000006B;
assign Y[4'b0001] [44] = 64'h000000000000042B;
assign u[4'b0001] [44] = 64'h000000000000082B;
assign v[4'b0001] [44] = 64'h0000000000000C2B;
assign X[4'b0001] [45] = 64'h000000000000006C;
assign Y[4'b0001] [45] = 64'h000000000000042C;
assign u[4'b0001] [45] = 64'h000000000000082C;
assign v[4'b0001] [45] = 64'h0000000000000C2C;
assign X[4'b0001] [46] = 64'h000000000000006D;
assign Y[4'b0001] [46] = 64'h000000000000042D;
assign u[4'b0001] [46] = 64'h000000000000082D;
assign v[4'b0001] [46] = 64'h0000000000000C2D;
assign X[4'b0001] [47] = 64'h000000000000006E;
assign Y[4'b0001] [47] = 64'h000000000000042E;
assign u[4'b0001] [47] = 64'h000000000000082E;
assign v[4'b0001] [47] = 64'h0000000000000C2E;
assign X[4'b0001] [48] = 64'h000000000000006F;
assign Y[4'b0001] [48] = 64'h000000000000042F;
assign u[4'b0001] [48] = 64'h000000000000082F;
assign v[4'b0001] [48] = 64'h0000000000000C2F;
assign X[4'b0001] [49] = 64'h0000000000000070;
assign Y[4'b0001] [49] = 64'h0000000000000430;
assign u[4'b0001] [49] = 64'h0000000000000830;
assign v[4'b0001] [49] = 64'h0000000000000C30;
assign X[4'b0001] [50] = 64'h0000000000000071;
assign Y[4'b0001] [50] = 64'h0000000000000431;
assign u[4'b0001] [50] = 64'h0000000000000831;
assign v[4'b0001] [50] = 64'h0000000000000C31;
assign X[4'b0001] [51] = 64'h0000000000000072;
assign Y[4'b0001] [51] = 64'h0000000000000432;
assign u[4'b0001] [51] = 64'h0000000000000832;
assign v[4'b0001] [51] = 64'h0000000000000C32;
assign X[4'b0001] [52] = 64'h0000000000000073;
assign Y[4'b0001] [52] = 64'h0000000000000433;
assign u[4'b0001] [52] = 64'h0000000000000833;
assign v[4'b0001] [52] = 64'h0000000000000C33;
assign X[4'b0001] [53] = 64'h0000000000000074;
assign Y[4'b0001] [53] = 64'h0000000000000434;
assign u[4'b0001] [53] = 64'h0000000000000834;
assign v[4'b0001] [53] = 64'h0000000000000C34;
assign X[4'b0001] [54] = 64'h0000000000000075;
assign Y[4'b0001] [54] = 64'h0000000000000435;
assign u[4'b0001] [54] = 64'h0000000000000835;
assign v[4'b0001] [54] = 64'h0000000000000C35;
assign X[4'b0001] [55] = 64'h0000000000000076;
assign Y[4'b0001] [55] = 64'h0000000000000436;
assign u[4'b0001] [55] = 64'h0000000000000836;
assign v[4'b0001] [55] = 64'h0000000000000C36;
assign X[4'b0001] [56] = 64'h0000000000000077;
assign Y[4'b0001] [56] = 64'h0000000000000437;
assign u[4'b0001] [56] = 64'h0000000000000837;
assign v[4'b0001] [56] = 64'h0000000000000C37;
assign X[4'b0001] [57] = 64'h0000000000000078;
assign Y[4'b0001] [57] = 64'h0000000000000438;
assign u[4'b0001] [57] = 64'h0000000000000838;
assign v[4'b0001] [57] = 64'h0000000000000C38;
assign X[4'b0001] [58] = 64'h0000000000000079;
assign Y[4'b0001] [58] = 64'h0000000000000439;
assign u[4'b0001] [58] = 64'h0000000000000839;
assign v[4'b0001] [58] = 64'h0000000000000C39;
assign X[4'b0001] [59] = 64'h000000000000007A;
assign Y[4'b0001] [59] = 64'h000000000000043A;
assign u[4'b0001] [59] = 64'h000000000000083A;
assign v[4'b0001] [59] = 64'h0000000000000C3A;
assign X[4'b0001] [60] = 64'h000000000000007B;
assign Y[4'b0001] [60] = 64'h000000000000043B;
assign u[4'b0001] [60] = 64'h000000000000083B;
assign v[4'b0001] [60] = 64'h0000000000000C3B;
assign X[4'b0001] [61] = 64'h000000000000007C;
assign Y[4'b0001] [61] = 64'h000000000000043C;
assign u[4'b0001] [61] = 64'h000000000000083C;
assign v[4'b0001] [61] = 64'h0000000000000C3C;
assign X[4'b0001] [62] = 64'h000000000000007D;
assign Y[4'b0001] [62] = 64'h000000000000043D;
assign u[4'b0001] [62] = 64'h000000000000083D;
assign v[4'b0001] [62] = 64'h0000000000000C3D;
assign X[4'b0001] [63] = 64'h000000000000007E;
assign Y[4'b0001] [63] = 64'h000000000000043E;
assign u[4'b0001] [63] = 64'h000000000000083E;
assign v[4'b0001] [63] = 64'h0000000000000C3E;
assign X[4'b0001] [64] = 64'h000000000000007F;
assign Y[4'b0001] [64] = 64'h000000000000043F;
assign u[4'b0001] [64] = 64'h000000000000083F;
assign v[4'b0001] [64] = 64'h0000000000000C3F;
assign X[4'b0010] [01] = 64'h0000000000000080;
assign Y[4'b0010] [01] = 64'h0000000000000440;
assign u[4'b0010] [01] = 64'h0000000000000840;
assign v[4'b0010] [01] = 64'h0000000000000C40;
assign X[4'b0010] [02] = 64'h0000000000000081;
assign Y[4'b0010] [02] = 64'h0000000000000441;
assign u[4'b0010] [02] = 64'h0000000000000841;
assign v[4'b0010] [02] = 64'h0000000000000C41;
assign X[4'b0010] [03] = 64'h0000000000000082;
assign Y[4'b0010] [03] = 64'h0000000000000442;
assign u[4'b0010] [03] = 64'h0000000000000842;
assign v[4'b0010] [03] = 64'h0000000000000C42;
assign X[4'b0010] [04] = 64'h0000000000000083;
assign Y[4'b0010] [04] = 64'h0000000000000443;
assign u[4'b0010] [04] = 64'h0000000000000843;
assign v[4'b0010] [04] = 64'h0000000000000C43;
assign X[4'b0010] [05] = 64'h0000000000000084;
assign Y[4'b0010] [05] = 64'h0000000000000444;
assign u[4'b0010] [05] = 64'h0000000000000844;
assign v[4'b0010] [05] = 64'h0000000000000C44;
assign X[4'b0010] [06] = 64'h0000000000000085;
assign Y[4'b0010] [06] = 64'h0000000000000445;
assign u[4'b0010] [06] = 64'h0000000000000845;
assign v[4'b0010] [06] = 64'h0000000000000C45;
assign X[4'b0010] [07] = 64'h0000000000000086;
assign Y[4'b0010] [07] = 64'h0000000000000446;
assign u[4'b0010] [07] = 64'h0000000000000846;
assign v[4'b0010] [07] = 64'h0000000000000C46;
assign X[4'b0010] [08] = 64'h0000000000000087;
assign Y[4'b0010] [08] = 64'h0000000000000447;
assign u[4'b0010] [08] = 64'h0000000000000847;
assign v[4'b0010] [08] = 64'h0000000000000C47;
assign X[4'b0010] [09] = 64'h0000000000000088;
assign Y[4'b0010] [09] = 64'h0000000000000448;
assign u[4'b0010] [09] = 64'h0000000000000848;
assign v[4'b0010] [09] = 64'h0000000000000C48;
assign X[4'b0010] [10] = 64'h0000000000000089;
assign Y[4'b0010] [10] = 64'h0000000000000449;
assign u[4'b0010] [10] = 64'h0000000000000849;
assign v[4'b0010] [10] = 64'h0000000000000C49;
assign X[4'b0010] [11] = 64'h000000000000008A;
assign Y[4'b0010] [11] = 64'h000000000000044A;
assign u[4'b0010] [11] = 64'h000000000000084A;
assign v[4'b0010] [11] = 64'h0000000000000C4A;
assign X[4'b0010] [12] = 64'h000000000000008B;
assign Y[4'b0010] [12] = 64'h000000000000044B;
assign u[4'b0010] [12] = 64'h000000000000084B;
assign v[4'b0010] [12] = 64'h0000000000000C4B;
assign X[4'b0010] [13] = 64'h000000000000008C;
assign Y[4'b0010] [13] = 64'h000000000000044C;
assign u[4'b0010] [13] = 64'h000000000000084C;
assign v[4'b0010] [13] = 64'h0000000000000C4C;
assign X[4'b0010] [14] = 64'h000000000000008D;
assign Y[4'b0010] [14] = 64'h000000000000044D;
assign u[4'b0010] [14] = 64'h000000000000084D;
assign v[4'b0010] [14] = 64'h0000000000000C4D;
assign X[4'b0010] [15] = 64'h000000000000008E;
assign Y[4'b0010] [15] = 64'h000000000000044E;
assign u[4'b0010] [15] = 64'h000000000000084E;
assign v[4'b0010] [15] = 64'h0000000000000C4E;
assign X[4'b0010] [16] = 64'h000000000000008F;
assign Y[4'b0010] [16] = 64'h000000000000044F;
assign u[4'b0010] [16] = 64'h000000000000084F;
assign v[4'b0010] [16] = 64'h0000000000000C4F;
assign X[4'b0010] [17] = 64'h0000000000000090;
assign Y[4'b0010] [17] = 64'h0000000000000450;
assign u[4'b0010] [17] = 64'h0000000000000850;
assign v[4'b0010] [17] = 64'h0000000000000C50;
assign X[4'b0010] [18] = 64'h0000000000000091;
assign Y[4'b0010] [18] = 64'h0000000000000451;
assign u[4'b0010] [18] = 64'h0000000000000851;
assign v[4'b0010] [18] = 64'h0000000000000C51;
assign X[4'b0010] [19] = 64'h0000000000000092;
assign Y[4'b0010] [19] = 64'h0000000000000452;
assign u[4'b0010] [19] = 64'h0000000000000852;
assign v[4'b0010] [19] = 64'h0000000000000C52;
assign X[4'b0010] [20] = 64'h0000000000000093;
assign Y[4'b0010] [20] = 64'h0000000000000453;
assign u[4'b0010] [20] = 64'h0000000000000853;
assign v[4'b0010] [20] = 64'h0000000000000C53;
assign X[4'b0010] [21] = 64'h0000000000000094;
assign Y[4'b0010] [21] = 64'h0000000000000454;
assign u[4'b0010] [21] = 64'h0000000000000854;
assign v[4'b0010] [21] = 64'h0000000000000C54;
assign X[4'b0010] [22] = 64'h0000000000000095;
assign Y[4'b0010] [22] = 64'h0000000000000455;
assign u[4'b0010] [22] = 64'h0000000000000855;
assign v[4'b0010] [22] = 64'h0000000000000C55;
assign X[4'b0010] [23] = 64'h0000000000000096;
assign Y[4'b0010] [23] = 64'h0000000000000456;
assign u[4'b0010] [23] = 64'h0000000000000856;
assign v[4'b0010] [23] = 64'h0000000000000C56;
assign X[4'b0010] [24] = 64'h0000000000000097;
assign Y[4'b0010] [24] = 64'h0000000000000457;
assign u[4'b0010] [24] = 64'h0000000000000857;
assign v[4'b0010] [24] = 64'h0000000000000C57;
assign X[4'b0010] [25] = 64'h0000000000000098;
assign Y[4'b0010] [25] = 64'h0000000000000458;
assign u[4'b0010] [25] = 64'h0000000000000858;
assign v[4'b0010] [25] = 64'h0000000000000C58;
assign X[4'b0010] [26] = 64'h0000000000000099;
assign Y[4'b0010] [26] = 64'h0000000000000459;
assign u[4'b0010] [26] = 64'h0000000000000859;
assign v[4'b0010] [26] = 64'h0000000000000C59;
assign X[4'b0010] [27] = 64'h000000000000009A;
assign Y[4'b0010] [27] = 64'h000000000000045A;
assign u[4'b0010] [27] = 64'h000000000000085A;
assign v[4'b0010] [27] = 64'h0000000000000C5A;
assign X[4'b0010] [28] = 64'h000000000000009B;
assign Y[4'b0010] [28] = 64'h000000000000045B;
assign u[4'b0010] [28] = 64'h000000000000085B;
assign v[4'b0010] [28] = 64'h0000000000000C5B;
assign X[4'b0010] [29] = 64'h000000000000009C;
assign Y[4'b0010] [29] = 64'h000000000000045C;
assign u[4'b0010] [29] = 64'h000000000000085C;
assign v[4'b0010] [29] = 64'h0000000000000C5C;
assign X[4'b0010] [30] = 64'h000000000000009D;
assign Y[4'b0010] [30] = 64'h000000000000045D;
assign u[4'b0010] [30] = 64'h000000000000085D;
assign v[4'b0010] [30] = 64'h0000000000000C5D;
assign X[4'b0010] [31] = 64'h000000000000009E;
assign Y[4'b0010] [31] = 64'h000000000000045E;
assign u[4'b0010] [31] = 64'h000000000000085E;
assign v[4'b0010] [31] = 64'h0000000000000C5E;
assign X[4'b0010] [32] = 64'h000000000000009F;
assign Y[4'b0010] [32] = 64'h000000000000045F;
assign u[4'b0010] [32] = 64'h000000000000085F;
assign v[4'b0010] [32] = 64'h0000000000000C5F;
assign X[4'b0010] [33] = 64'h00000000000000A0;
assign Y[4'b0010] [33] = 64'h0000000000000460;
assign u[4'b0010] [33] = 64'h0000000000000860;
assign v[4'b0010] [33] = 64'h0000000000000C60;
assign X[4'b0010] [34] = 64'h00000000000000A1;
assign Y[4'b0010] [34] = 64'h0000000000000461;
assign u[4'b0010] [34] = 64'h0000000000000861;
assign v[4'b0010] [34] = 64'h0000000000000C61;
assign X[4'b0010] [35] = 64'h00000000000000A2;
assign Y[4'b0010] [35] = 64'h0000000000000462;
assign u[4'b0010] [35] = 64'h0000000000000862;
assign v[4'b0010] [35] = 64'h0000000000000C62;
assign X[4'b0010] [36] = 64'h00000000000000A3;
assign Y[4'b0010] [36] = 64'h0000000000000463;
assign u[4'b0010] [36] = 64'h0000000000000863;
assign v[4'b0010] [36] = 64'h0000000000000C63;
assign X[4'b0010] [37] = 64'h00000000000000A4;
assign Y[4'b0010] [37] = 64'h0000000000000464;
assign u[4'b0010] [37] = 64'h0000000000000864;
assign v[4'b0010] [37] = 64'h0000000000000C64;
assign X[4'b0010] [38] = 64'h00000000000000A5;
assign Y[4'b0010] [38] = 64'h0000000000000465;
assign u[4'b0010] [38] = 64'h0000000000000865;
assign v[4'b0010] [38] = 64'h0000000000000C65;
assign X[4'b0010] [39] = 64'h00000000000000A6;
assign Y[4'b0010] [39] = 64'h0000000000000466;
assign u[4'b0010] [39] = 64'h0000000000000866;
assign v[4'b0010] [39] = 64'h0000000000000C66;
assign X[4'b0010] [40] = 64'h00000000000000A7;
assign Y[4'b0010] [40] = 64'h0000000000000467;
assign u[4'b0010] [40] = 64'h0000000000000867;
assign v[4'b0010] [40] = 64'h0000000000000C67;
assign X[4'b0010] [41] = 64'h00000000000000A8;
assign Y[4'b0010] [41] = 64'h0000000000000468;
assign u[4'b0010] [41] = 64'h0000000000000868;
assign v[4'b0010] [41] = 64'h0000000000000C68;
assign X[4'b0010] [42] = 64'h00000000000000A9;
assign Y[4'b0010] [42] = 64'h0000000000000469;
assign u[4'b0010] [42] = 64'h0000000000000869;
assign v[4'b0010] [42] = 64'h0000000000000C69;
assign X[4'b0010] [43] = 64'h00000000000000AA;
assign Y[4'b0010] [43] = 64'h000000000000046A;
assign u[4'b0010] [43] = 64'h000000000000086A;
assign v[4'b0010] [43] = 64'h0000000000000C6A;
assign X[4'b0010] [44] = 64'h00000000000000AB;
assign Y[4'b0010] [44] = 64'h000000000000046B;
assign u[4'b0010] [44] = 64'h000000000000086B;
assign v[4'b0010] [44] = 64'h0000000000000C6B;
assign X[4'b0010] [45] = 64'h00000000000000AC;
assign Y[4'b0010] [45] = 64'h000000000000046C;
assign u[4'b0010] [45] = 64'h000000000000086C;
assign v[4'b0010] [45] = 64'h0000000000000C6C;
assign X[4'b0010] [46] = 64'h00000000000000AD;
assign Y[4'b0010] [46] = 64'h000000000000046D;
assign u[4'b0010] [46] = 64'h000000000000086D;
assign v[4'b0010] [46] = 64'h0000000000000C6D;
assign X[4'b0010] [47] = 64'h00000000000000AE;
assign Y[4'b0010] [47] = 64'h000000000000046E;
assign u[4'b0010] [47] = 64'h000000000000086E;
assign v[4'b0010] [47] = 64'h0000000000000C6E;
assign X[4'b0010] [48] = 64'h00000000000000AF;
assign Y[4'b0010] [48] = 64'h000000000000046F;
assign u[4'b0010] [48] = 64'h000000000000086F;
assign v[4'b0010] [48] = 64'h0000000000000C6F;
assign X[4'b0010] [49] = 64'h00000000000000B0;
assign Y[4'b0010] [49] = 64'h0000000000000470;
assign u[4'b0010] [49] = 64'h0000000000000870;
assign v[4'b0010] [49] = 64'h0000000000000C70;
assign X[4'b0010] [50] = 64'h00000000000000B1;
assign Y[4'b0010] [50] = 64'h0000000000000471;
assign u[4'b0010] [50] = 64'h0000000000000871;
assign v[4'b0010] [50] = 64'h0000000000000C71;
assign X[4'b0010] [51] = 64'h00000000000000B2;
assign Y[4'b0010] [51] = 64'h0000000000000472;
assign u[4'b0010] [51] = 64'h0000000000000872;
assign v[4'b0010] [51] = 64'h0000000000000C72;
assign X[4'b0010] [52] = 64'h00000000000000B3;
assign Y[4'b0010] [52] = 64'h0000000000000473;
assign u[4'b0010] [52] = 64'h0000000000000873;
assign v[4'b0010] [52] = 64'h0000000000000C73;
assign X[4'b0010] [53] = 64'h00000000000000B4;
assign Y[4'b0010] [53] = 64'h0000000000000474;
assign u[4'b0010] [53] = 64'h0000000000000874;
assign v[4'b0010] [53] = 64'h0000000000000C74;
assign X[4'b0010] [54] = 64'h00000000000000B5;
assign Y[4'b0010] [54] = 64'h0000000000000475;
assign u[4'b0010] [54] = 64'h0000000000000875;
assign v[4'b0010] [54] = 64'h0000000000000C75;
assign X[4'b0010] [55] = 64'h00000000000000B6;
assign Y[4'b0010] [55] = 64'h0000000000000476;
assign u[4'b0010] [55] = 64'h0000000000000876;
assign v[4'b0010] [55] = 64'h0000000000000C76;
assign X[4'b0010] [56] = 64'h00000000000000B7;
assign Y[4'b0010] [56] = 64'h0000000000000477;
assign u[4'b0010] [56] = 64'h0000000000000877;
assign v[4'b0010] [56] = 64'h0000000000000C77;
assign X[4'b0010] [57] = 64'h00000000000000B8;
assign Y[4'b0010] [57] = 64'h0000000000000478;
assign u[4'b0010] [57] = 64'h0000000000000878;
assign v[4'b0010] [57] = 64'h0000000000000C78;
assign X[4'b0010] [58] = 64'h00000000000000B9;
assign Y[4'b0010] [58] = 64'h0000000000000479;
assign u[4'b0010] [58] = 64'h0000000000000879;
assign v[4'b0010] [58] = 64'h0000000000000C79;
assign X[4'b0010] [59] = 64'h00000000000000BA;
assign Y[4'b0010] [59] = 64'h000000000000047A;
assign u[4'b0010] [59] = 64'h000000000000087A;
assign v[4'b0010] [59] = 64'h0000000000000C7A;
assign X[4'b0010] [60] = 64'h00000000000000BB;
assign Y[4'b0010] [60] = 64'h000000000000047B;
assign u[4'b0010] [60] = 64'h000000000000087B;
assign v[4'b0010] [60] = 64'h0000000000000C7B;
assign X[4'b0010] [61] = 64'h00000000000000BC;
assign Y[4'b0010] [61] = 64'h000000000000047C;
assign u[4'b0010] [61] = 64'h000000000000087C;
assign v[4'b0010] [61] = 64'h0000000000000C7C;
assign X[4'b0010] [62] = 64'h00000000000000BD;
assign Y[4'b0010] [62] = 64'h000000000000047D;
assign u[4'b0010] [62] = 64'h000000000000087D;
assign v[4'b0010] [62] = 64'h0000000000000C7D;
assign X[4'b0010] [63] = 64'h00000000000000BE;
assign Y[4'b0010] [63] = 64'h000000000000047E;
assign u[4'b0010] [63] = 64'h000000000000087E;
assign v[4'b0010] [63] = 64'h0000000000000C7E;
assign X[4'b0010] [64] = 64'h00000000000000BF;
assign Y[4'b0010] [64] = 64'h000000000000047F;
assign u[4'b0010] [64] = 64'h000000000000087F;
assign v[4'b0010] [64] = 64'h0000000000000C7F;
assign X[4'b0011] [01] = 64'h00000000000000C0;
assign Y[4'b0011] [01] = 64'h0000000000000480;
assign u[4'b0011] [01] = 64'h0000000000000880;
assign v[4'b0011] [01] = 64'h0000000000000C80;
assign X[4'b0011] [02] = 64'h00000000000000C1;
assign Y[4'b0011] [02] = 64'h0000000000000481;
assign u[4'b0011] [02] = 64'h0000000000000881;
assign v[4'b0011] [02] = 64'h0000000000000C81;
assign X[4'b0011] [03] = 64'h00000000000000C2;
assign Y[4'b0011] [03] = 64'h0000000000000482;
assign u[4'b0011] [03] = 64'h0000000000000882;
assign v[4'b0011] [03] = 64'h0000000000000C82;
assign X[4'b0011] [04] = 64'h00000000000000C3;
assign Y[4'b0011] [04] = 64'h0000000000000483;
assign u[4'b0011] [04] = 64'h0000000000000883;
assign v[4'b0011] [04] = 64'h0000000000000C83;
assign X[4'b0011] [05] = 64'h00000000000000C4;
assign Y[4'b0011] [05] = 64'h0000000000000484;
assign u[4'b0011] [05] = 64'h0000000000000884;
assign v[4'b0011] [05] = 64'h0000000000000C84;
assign X[4'b0011] [06] = 64'h00000000000000C5;
assign Y[4'b0011] [06] = 64'h0000000000000485;
assign u[4'b0011] [06] = 64'h0000000000000885;
assign v[4'b0011] [06] = 64'h0000000000000C85;
assign X[4'b0011] [07] = 64'h00000000000000C6;
assign Y[4'b0011] [07] = 64'h0000000000000486;
assign u[4'b0011] [07] = 64'h0000000000000886;
assign v[4'b0011] [07] = 64'h0000000000000C86;
assign X[4'b0011] [08] = 64'h00000000000000C7;
assign Y[4'b0011] [08] = 64'h0000000000000487;
assign u[4'b0011] [08] = 64'h0000000000000887;
assign v[4'b0011] [08] = 64'h0000000000000C87;
assign X[4'b0011] [09] = 64'h00000000000000C8;
assign Y[4'b0011] [09] = 64'h0000000000000488;
assign u[4'b0011] [09] = 64'h0000000000000888;
assign v[4'b0011] [09] = 64'h0000000000000C88;
assign X[4'b0011] [10] = 64'h00000000000000C9;
assign Y[4'b0011] [10] = 64'h0000000000000489;
assign u[4'b0011] [10] = 64'h0000000000000889;
assign v[4'b0011] [10] = 64'h0000000000000C89;
assign X[4'b0011] [11] = 64'h00000000000000CA;
assign Y[4'b0011] [11] = 64'h000000000000048A;
assign u[4'b0011] [11] = 64'h000000000000088A;
assign v[4'b0011] [11] = 64'h0000000000000C8A;
assign X[4'b0011] [12] = 64'h00000000000000CB;
assign Y[4'b0011] [12] = 64'h000000000000048B;
assign u[4'b0011] [12] = 64'h000000000000088B;
assign v[4'b0011] [12] = 64'h0000000000000C8B;
assign X[4'b0011] [13] = 64'h00000000000000CC;
assign Y[4'b0011] [13] = 64'h000000000000048C;
assign u[4'b0011] [13] = 64'h000000000000088C;
assign v[4'b0011] [13] = 64'h0000000000000C8C;
assign X[4'b0011] [14] = 64'h00000000000000CD;
assign Y[4'b0011] [14] = 64'h000000000000048D;
assign u[4'b0011] [14] = 64'h000000000000088D;
assign v[4'b0011] [14] = 64'h0000000000000C8D;
assign X[4'b0011] [15] = 64'h00000000000000CE;
assign Y[4'b0011] [15] = 64'h000000000000048E;
assign u[4'b0011] [15] = 64'h000000000000088E;
assign v[4'b0011] [15] = 64'h0000000000000C8E;
assign X[4'b0011] [16] = 64'h00000000000000CF;
assign Y[4'b0011] [16] = 64'h000000000000048F;
assign u[4'b0011] [16] = 64'h000000000000088F;
assign v[4'b0011] [16] = 64'h0000000000000C8F;
assign X[4'b0011] [17] = 64'h00000000000000D0;
assign Y[4'b0011] [17] = 64'h0000000000000490;
assign u[4'b0011] [17] = 64'h0000000000000890;
assign v[4'b0011] [17] = 64'h0000000000000C90;
assign X[4'b0011] [18] = 64'h00000000000000D1;
assign Y[4'b0011] [18] = 64'h0000000000000491;
assign u[4'b0011] [18] = 64'h0000000000000891;
assign v[4'b0011] [18] = 64'h0000000000000C91;
assign X[4'b0011] [19] = 64'h00000000000000D2;
assign Y[4'b0011] [19] = 64'h0000000000000492;
assign u[4'b0011] [19] = 64'h0000000000000892;
assign v[4'b0011] [19] = 64'h0000000000000C92;
assign X[4'b0011] [20] = 64'h00000000000000D3;
assign Y[4'b0011] [20] = 64'h0000000000000493;
assign u[4'b0011] [20] = 64'h0000000000000893;
assign v[4'b0011] [20] = 64'h0000000000000C93;
assign X[4'b0011] [21] = 64'h00000000000000D4;
assign Y[4'b0011] [21] = 64'h0000000000000494;
assign u[4'b0011] [21] = 64'h0000000000000894;
assign v[4'b0011] [21] = 64'h0000000000000C94;
assign X[4'b0011] [22] = 64'h00000000000000D5;
assign Y[4'b0011] [22] = 64'h0000000000000495;
assign u[4'b0011] [22] = 64'h0000000000000895;
assign v[4'b0011] [22] = 64'h0000000000000C95;
assign X[4'b0011] [23] = 64'h00000000000000D6;
assign Y[4'b0011] [23] = 64'h0000000000000496;
assign u[4'b0011] [23] = 64'h0000000000000896;
assign v[4'b0011] [23] = 64'h0000000000000C96;
assign X[4'b0011] [24] = 64'h00000000000000D7;
assign Y[4'b0011] [24] = 64'h0000000000000497;
assign u[4'b0011] [24] = 64'h0000000000000897;
assign v[4'b0011] [24] = 64'h0000000000000C97;
assign X[4'b0011] [25] = 64'h00000000000000D8;
assign Y[4'b0011] [25] = 64'h0000000000000498;
assign u[4'b0011] [25] = 64'h0000000000000898;
assign v[4'b0011] [25] = 64'h0000000000000C98;
assign X[4'b0011] [26] = 64'h00000000000000D9;
assign Y[4'b0011] [26] = 64'h0000000000000499;
assign u[4'b0011] [26] = 64'h0000000000000899;
assign v[4'b0011] [26] = 64'h0000000000000C99;
assign X[4'b0011] [27] = 64'h00000000000000DA;
assign Y[4'b0011] [27] = 64'h000000000000049A;
assign u[4'b0011] [27] = 64'h000000000000089A;
assign v[4'b0011] [27] = 64'h0000000000000C9A;
assign X[4'b0011] [28] = 64'h00000000000000DB;
assign Y[4'b0011] [28] = 64'h000000000000049B;
assign u[4'b0011] [28] = 64'h000000000000089B;
assign v[4'b0011] [28] = 64'h0000000000000C9B;
assign X[4'b0011] [29] = 64'h00000000000000DC;
assign Y[4'b0011] [29] = 64'h000000000000049C;
assign u[4'b0011] [29] = 64'h000000000000089C;
assign v[4'b0011] [29] = 64'h0000000000000C9C;
assign X[4'b0011] [30] = 64'h00000000000000DD;
assign Y[4'b0011] [30] = 64'h000000000000049D;
assign u[4'b0011] [30] = 64'h000000000000089D;
assign v[4'b0011] [30] = 64'h0000000000000C9D;
assign X[4'b0011] [31] = 64'h00000000000000DE;
assign Y[4'b0011] [31] = 64'h000000000000049E;
assign u[4'b0011] [31] = 64'h000000000000089E;
assign v[4'b0011] [31] = 64'h0000000000000C9E;
assign X[4'b0011] [32] = 64'h00000000000000DF;
assign Y[4'b0011] [32] = 64'h000000000000049F;
assign u[4'b0011] [32] = 64'h000000000000089F;
assign v[4'b0011] [32] = 64'h0000000000000C9F;
assign X[4'b0011] [33] = 64'h00000000000000E0;
assign Y[4'b0011] [33] = 64'h00000000000004A0;
assign u[4'b0011] [33] = 64'h00000000000008A0;
assign v[4'b0011] [33] = 64'h0000000000000CA0;
assign X[4'b0011] [34] = 64'h00000000000000E1;
assign Y[4'b0011] [34] = 64'h00000000000004A1;
assign u[4'b0011] [34] = 64'h00000000000008A1;
assign v[4'b0011] [34] = 64'h0000000000000CA1;
assign X[4'b0011] [35] = 64'h00000000000000E2;
assign Y[4'b0011] [35] = 64'h00000000000004A2;
assign u[4'b0011] [35] = 64'h00000000000008A2;
assign v[4'b0011] [35] = 64'h0000000000000CA2;
assign X[4'b0011] [36] = 64'h00000000000000E3;
assign Y[4'b0011] [36] = 64'h00000000000004A3;
assign u[4'b0011] [36] = 64'h00000000000008A3;
assign v[4'b0011] [36] = 64'h0000000000000CA3;
assign X[4'b0011] [37] = 64'h00000000000000E4;
assign Y[4'b0011] [37] = 64'h00000000000004A4;
assign u[4'b0011] [37] = 64'h00000000000008A4;
assign v[4'b0011] [37] = 64'h0000000000000CA4;
assign X[4'b0011] [38] = 64'h00000000000000E5;
assign Y[4'b0011] [38] = 64'h00000000000004A5;
assign u[4'b0011] [38] = 64'h00000000000008A5;
assign v[4'b0011] [38] = 64'h0000000000000CA5;
assign X[4'b0011] [39] = 64'h00000000000000E6;
assign Y[4'b0011] [39] = 64'h00000000000004A6;
assign u[4'b0011] [39] = 64'h00000000000008A6;
assign v[4'b0011] [39] = 64'h0000000000000CA6;
assign X[4'b0011] [40] = 64'h00000000000000E7;
assign Y[4'b0011] [40] = 64'h00000000000004A7;
assign u[4'b0011] [40] = 64'h00000000000008A7;
assign v[4'b0011] [40] = 64'h0000000000000CA7;
assign X[4'b0011] [41] = 64'h00000000000000E8;
assign Y[4'b0011] [41] = 64'h00000000000004A8;
assign u[4'b0011] [41] = 64'h00000000000008A8;
assign v[4'b0011] [41] = 64'h0000000000000CA8;
assign X[4'b0011] [42] = 64'h00000000000000E9;
assign Y[4'b0011] [42] = 64'h00000000000004A9;
assign u[4'b0011] [42] = 64'h00000000000008A9;
assign v[4'b0011] [42] = 64'h0000000000000CA9;
assign X[4'b0011] [43] = 64'h00000000000000EA;
assign Y[4'b0011] [43] = 64'h00000000000004AA;
assign u[4'b0011] [43] = 64'h00000000000008AA;
assign v[4'b0011] [43] = 64'h0000000000000CAA;
assign X[4'b0011] [44] = 64'h00000000000000EB;
assign Y[4'b0011] [44] = 64'h00000000000004AB;
assign u[4'b0011] [44] = 64'h00000000000008AB;
assign v[4'b0011] [44] = 64'h0000000000000CAB;
assign X[4'b0011] [45] = 64'h00000000000000EC;
assign Y[4'b0011] [45] = 64'h00000000000004AC;
assign u[4'b0011] [45] = 64'h00000000000008AC;
assign v[4'b0011] [45] = 64'h0000000000000CAC;
assign X[4'b0011] [46] = 64'h00000000000000ED;
assign Y[4'b0011] [46] = 64'h00000000000004AD;
assign u[4'b0011] [46] = 64'h00000000000008AD;
assign v[4'b0011] [46] = 64'h0000000000000CAD;
assign X[4'b0011] [47] = 64'h00000000000000EE;
assign Y[4'b0011] [47] = 64'h00000000000004AE;
assign u[4'b0011] [47] = 64'h00000000000008AE;
assign v[4'b0011] [47] = 64'h0000000000000CAE;
assign X[4'b0011] [48] = 64'h00000000000000EF;
assign Y[4'b0011] [48] = 64'h00000000000004AF;
assign u[4'b0011] [48] = 64'h00000000000008AF;
assign v[4'b0011] [48] = 64'h0000000000000CAF;
assign X[4'b0011] [49] = 64'h00000000000000F0;
assign Y[4'b0011] [49] = 64'h00000000000004B0;
assign u[4'b0011] [49] = 64'h00000000000008B0;
assign v[4'b0011] [49] = 64'h0000000000000CB0;
assign X[4'b0011] [50] = 64'h00000000000000F1;
assign Y[4'b0011] [50] = 64'h00000000000004B1;
assign u[4'b0011] [50] = 64'h00000000000008B1;
assign v[4'b0011] [50] = 64'h0000000000000CB1;
assign X[4'b0011] [51] = 64'h00000000000000F2;
assign Y[4'b0011] [51] = 64'h00000000000004B2;
assign u[4'b0011] [51] = 64'h00000000000008B2;
assign v[4'b0011] [51] = 64'h0000000000000CB2;
assign X[4'b0011] [52] = 64'h00000000000000F3;
assign Y[4'b0011] [52] = 64'h00000000000004B3;
assign u[4'b0011] [52] = 64'h00000000000008B3;
assign v[4'b0011] [52] = 64'h0000000000000CB3;
assign X[4'b0011] [53] = 64'h00000000000000F4;
assign Y[4'b0011] [53] = 64'h00000000000004B4;
assign u[4'b0011] [53] = 64'h00000000000008B4;
assign v[4'b0011] [53] = 64'h0000000000000CB4;
assign X[4'b0011] [54] = 64'h00000000000000F5;
assign Y[4'b0011] [54] = 64'h00000000000004B5;
assign u[4'b0011] [54] = 64'h00000000000008B5;
assign v[4'b0011] [54] = 64'h0000000000000CB5;
assign X[4'b0011] [55] = 64'h00000000000000F6;
assign Y[4'b0011] [55] = 64'h00000000000004B6;
assign u[4'b0011] [55] = 64'h00000000000008B6;
assign v[4'b0011] [55] = 64'h0000000000000CB6;
assign X[4'b0011] [56] = 64'h00000000000000F7;
assign Y[4'b0011] [56] = 64'h00000000000004B7;
assign u[4'b0011] [56] = 64'h00000000000008B7;
assign v[4'b0011] [56] = 64'h0000000000000CB7;
assign X[4'b0011] [57] = 64'h00000000000000F8;
assign Y[4'b0011] [57] = 64'h00000000000004B8;
assign u[4'b0011] [57] = 64'h00000000000008B8;
assign v[4'b0011] [57] = 64'h0000000000000CB8;
assign X[4'b0011] [58] = 64'h00000000000000F9;
assign Y[4'b0011] [58] = 64'h00000000000004B9;
assign u[4'b0011] [58] = 64'h00000000000008B9;
assign v[4'b0011] [58] = 64'h0000000000000CB9;
assign X[4'b0011] [59] = 64'h00000000000000FA;
assign Y[4'b0011] [59] = 64'h00000000000004BA;
assign u[4'b0011] [59] = 64'h00000000000008BA;
assign v[4'b0011] [59] = 64'h0000000000000CBA;
assign X[4'b0011] [60] = 64'h00000000000000FB;
assign Y[4'b0011] [60] = 64'h00000000000004BB;
assign u[4'b0011] [60] = 64'h00000000000008BB;
assign v[4'b0011] [60] = 64'h0000000000000CBB;
assign X[4'b0011] [61] = 64'h00000000000000FC;
assign Y[4'b0011] [61] = 64'h00000000000004BC;
assign u[4'b0011] [61] = 64'h00000000000008BC;
assign v[4'b0011] [61] = 64'h0000000000000CBC;
assign X[4'b0011] [62] = 64'h00000000000000FD;
assign Y[4'b0011] [62] = 64'h00000000000004BD;
assign u[4'b0011] [62] = 64'h00000000000008BD;
assign v[4'b0011] [62] = 64'h0000000000000CBD;
assign X[4'b0011] [63] = 64'h00000000000000FE;
assign Y[4'b0011] [63] = 64'h00000000000004BE;
assign u[4'b0011] [63] = 64'h00000000000008BE;
assign v[4'b0011] [63] = 64'h0000000000000CBE;
assign X[4'b0011] [64] = 64'h00000000000000FF;
assign Y[4'b0011] [64] = 64'h00000000000004BF;
assign u[4'b0011] [64] = 64'h00000000000008BF;
assign v[4'b0011] [64] = 64'h0000000000000CBF;
assign X[4'b0100] [01] = 64'h0000000000000100;
assign Y[4'b0100] [01] = 64'h00000000000004C0;
assign u[4'b0100] [01] = 64'h00000000000008C0;
assign v[4'b0100] [01] = 64'h0000000000000CC0;
assign X[4'b0100] [02] = 64'h0000000000000101;
assign Y[4'b0100] [02] = 64'h00000000000004C1;
assign u[4'b0100] [02] = 64'h00000000000008C1;
assign v[4'b0100] [02] = 64'h0000000000000CC1;
assign X[4'b0100] [03] = 64'h0000000000000102;
assign Y[4'b0100] [03] = 64'h00000000000004C2;
assign u[4'b0100] [03] = 64'h00000000000008C2;
assign v[4'b0100] [03] = 64'h0000000000000CC2;
assign X[4'b0100] [04] = 64'h0000000000000103;
assign Y[4'b0100] [04] = 64'h00000000000004C3;
assign u[4'b0100] [04] = 64'h00000000000008C3;
assign v[4'b0100] [04] = 64'h0000000000000CC3;
assign X[4'b0100] [05] = 64'h0000000000000104;
assign Y[4'b0100] [05] = 64'h00000000000004C4;
assign u[4'b0100] [05] = 64'h00000000000008C4;
assign v[4'b0100] [05] = 64'h0000000000000CC4;
assign X[4'b0100] [06] = 64'h0000000000000105;
assign Y[4'b0100] [06] = 64'h00000000000004C5;
assign u[4'b0100] [06] = 64'h00000000000008C5;
assign v[4'b0100] [06] = 64'h0000000000000CC5;
assign X[4'b0100] [07] = 64'h0000000000000106;
assign Y[4'b0100] [07] = 64'h00000000000004C6;
assign u[4'b0100] [07] = 64'h00000000000008C6;
assign v[4'b0100] [07] = 64'h0000000000000CC6;
assign X[4'b0100] [08] = 64'h0000000000000107;
assign Y[4'b0100] [08] = 64'h00000000000004C7;
assign u[4'b0100] [08] = 64'h00000000000008C7;
assign v[4'b0100] [08] = 64'h0000000000000CC7;
assign X[4'b0100] [09] = 64'h0000000000000108;
assign Y[4'b0100] [09] = 64'h00000000000004C8;
assign u[4'b0100] [09] = 64'h00000000000008C8;
assign v[4'b0100] [09] = 64'h0000000000000CC8;
assign X[4'b0100] [10] = 64'h0000000000000109;
assign Y[4'b0100] [10] = 64'h00000000000004C9;
assign u[4'b0100] [10] = 64'h00000000000008C9;
assign v[4'b0100] [10] = 64'h0000000000000CC9;
assign X[4'b0100] [11] = 64'h000000000000010A;
assign Y[4'b0100] [11] = 64'h00000000000004CA;
assign u[4'b0100] [11] = 64'h00000000000008CA;
assign v[4'b0100] [11] = 64'h0000000000000CCA;
assign X[4'b0100] [12] = 64'h000000000000010B;
assign Y[4'b0100] [12] = 64'h00000000000004CB;
assign u[4'b0100] [12] = 64'h00000000000008CB;
assign v[4'b0100] [12] = 64'h0000000000000CCB;
assign X[4'b0100] [13] = 64'h000000000000010C;
assign Y[4'b0100] [13] = 64'h00000000000004CC;
assign u[4'b0100] [13] = 64'h00000000000008CC;
assign v[4'b0100] [13] = 64'h0000000000000CCC;
assign X[4'b0100] [14] = 64'h000000000000010D;
assign Y[4'b0100] [14] = 64'h00000000000004CD;
assign u[4'b0100] [14] = 64'h00000000000008CD;
assign v[4'b0100] [14] = 64'h0000000000000CCD;
assign X[4'b0100] [15] = 64'h000000000000010E;
assign Y[4'b0100] [15] = 64'h00000000000004CE;
assign u[4'b0100] [15] = 64'h00000000000008CE;
assign v[4'b0100] [15] = 64'h0000000000000CCE;
assign X[4'b0100] [16] = 64'h000000000000010F;
assign Y[4'b0100] [16] = 64'h00000000000004CF;
assign u[4'b0100] [16] = 64'h00000000000008CF;
assign v[4'b0100] [16] = 64'h0000000000000CCF;
assign X[4'b0100] [17] = 64'h0000000000000110;
assign Y[4'b0100] [17] = 64'h00000000000004D0;
assign u[4'b0100] [17] = 64'h00000000000008D0;
assign v[4'b0100] [17] = 64'h0000000000000CD0;
assign X[4'b0100] [18] = 64'h0000000000000111;
assign Y[4'b0100] [18] = 64'h00000000000004D1;
assign u[4'b0100] [18] = 64'h00000000000008D1;
assign v[4'b0100] [18] = 64'h0000000000000CD1;
assign X[4'b0100] [19] = 64'h0000000000000112;
assign Y[4'b0100] [19] = 64'h00000000000004D2;
assign u[4'b0100] [19] = 64'h00000000000008D2;
assign v[4'b0100] [19] = 64'h0000000000000CD2;
assign X[4'b0100] [20] = 64'h0000000000000113;
assign Y[4'b0100] [20] = 64'h00000000000004D3;
assign u[4'b0100] [20] = 64'h00000000000008D3;
assign v[4'b0100] [20] = 64'h0000000000000CD3;
assign X[4'b0100] [21] = 64'h0000000000000114;
assign Y[4'b0100] [21] = 64'h00000000000004D4;
assign u[4'b0100] [21] = 64'h00000000000008D4;
assign v[4'b0100] [21] = 64'h0000000000000CD4;
assign X[4'b0100] [22] = 64'h0000000000000115;
assign Y[4'b0100] [22] = 64'h00000000000004D5;
assign u[4'b0100] [22] = 64'h00000000000008D5;
assign v[4'b0100] [22] = 64'h0000000000000CD5;
assign X[4'b0100] [23] = 64'h0000000000000116;
assign Y[4'b0100] [23] = 64'h00000000000004D6;
assign u[4'b0100] [23] = 64'h00000000000008D6;
assign v[4'b0100] [23] = 64'h0000000000000CD6;
assign X[4'b0100] [24] = 64'h0000000000000117;
assign Y[4'b0100] [24] = 64'h00000000000004D7;
assign u[4'b0100] [24] = 64'h00000000000008D7;
assign v[4'b0100] [24] = 64'h0000000000000CD7;
assign X[4'b0100] [25] = 64'h0000000000000118;
assign Y[4'b0100] [25] = 64'h00000000000004D8;
assign u[4'b0100] [25] = 64'h00000000000008D8;
assign v[4'b0100] [25] = 64'h0000000000000CD8;
assign X[4'b0100] [26] = 64'h0000000000000119;
assign Y[4'b0100] [26] = 64'h00000000000004D9;
assign u[4'b0100] [26] = 64'h00000000000008D9;
assign v[4'b0100] [26] = 64'h0000000000000CD9;
assign X[4'b0100] [27] = 64'h000000000000011A;
assign Y[4'b0100] [27] = 64'h00000000000004DA;
assign u[4'b0100] [27] = 64'h00000000000008DA;
assign v[4'b0100] [27] = 64'h0000000000000CDA;
assign X[4'b0100] [28] = 64'h000000000000011B;
assign Y[4'b0100] [28] = 64'h00000000000004DB;
assign u[4'b0100] [28] = 64'h00000000000008DB;
assign v[4'b0100] [28] = 64'h0000000000000CDB;
assign X[4'b0100] [29] = 64'h000000000000011C;
assign Y[4'b0100] [29] = 64'h00000000000004DC;
assign u[4'b0100] [29] = 64'h00000000000008DC;
assign v[4'b0100] [29] = 64'h0000000000000CDC;
assign X[4'b0100] [30] = 64'h000000000000011D;
assign Y[4'b0100] [30] = 64'h00000000000004DD;
assign u[4'b0100] [30] = 64'h00000000000008DD;
assign v[4'b0100] [30] = 64'h0000000000000CDD;
assign X[4'b0100] [31] = 64'h000000000000011E;
assign Y[4'b0100] [31] = 64'h00000000000004DE;
assign u[4'b0100] [31] = 64'h00000000000008DE;
assign v[4'b0100] [31] = 64'h0000000000000CDE;
assign X[4'b0100] [32] = 64'h000000000000011F;
assign Y[4'b0100] [32] = 64'h00000000000004DF;
assign u[4'b0100] [32] = 64'h00000000000008DF;
assign v[4'b0100] [32] = 64'h0000000000000CDF;
assign X[4'b0100] [33] = 64'h0000000000000120;
assign Y[4'b0100] [33] = 64'h00000000000004E0;
assign u[4'b0100] [33] = 64'h00000000000008E0;
assign v[4'b0100] [33] = 64'h0000000000000CE0;
assign X[4'b0100] [34] = 64'h0000000000000121;
assign Y[4'b0100] [34] = 64'h00000000000004E1;
assign u[4'b0100] [34] = 64'h00000000000008E1;
assign v[4'b0100] [34] = 64'h0000000000000CE1;
assign X[4'b0100] [35] = 64'h0000000000000122;
assign Y[4'b0100] [35] = 64'h00000000000004E2;
assign u[4'b0100] [35] = 64'h00000000000008E2;
assign v[4'b0100] [35] = 64'h0000000000000CE2;
assign X[4'b0100] [36] = 64'h0000000000000123;
assign Y[4'b0100] [36] = 64'h00000000000004E3;
assign u[4'b0100] [36] = 64'h00000000000008E3;
assign v[4'b0100] [36] = 64'h0000000000000CE3;
assign X[4'b0100] [37] = 64'h0000000000000124;
assign Y[4'b0100] [37] = 64'h00000000000004E4;
assign u[4'b0100] [37] = 64'h00000000000008E4;
assign v[4'b0100] [37] = 64'h0000000000000CE4;
assign X[4'b0100] [38] = 64'h0000000000000125;
assign Y[4'b0100] [38] = 64'h00000000000004E5;
assign u[4'b0100] [38] = 64'h00000000000008E5;
assign v[4'b0100] [38] = 64'h0000000000000CE5;
assign X[4'b0100] [39] = 64'h0000000000000126;
assign Y[4'b0100] [39] = 64'h00000000000004E6;
assign u[4'b0100] [39] = 64'h00000000000008E6;
assign v[4'b0100] [39] = 64'h0000000000000CE6;
assign X[4'b0100] [40] = 64'h0000000000000127;
assign Y[4'b0100] [40] = 64'h00000000000004E7;
assign u[4'b0100] [40] = 64'h00000000000008E7;
assign v[4'b0100] [40] = 64'h0000000000000CE7;
assign X[4'b0100] [41] = 64'h0000000000000128;
assign Y[4'b0100] [41] = 64'h00000000000004E8;
assign u[4'b0100] [41] = 64'h00000000000008E8;
assign v[4'b0100] [41] = 64'h0000000000000CE8;
assign X[4'b0100] [42] = 64'h0000000000000129;
assign Y[4'b0100] [42] = 64'h00000000000004E9;
assign u[4'b0100] [42] = 64'h00000000000008E9;
assign v[4'b0100] [42] = 64'h0000000000000CE9;
assign X[4'b0100] [43] = 64'h000000000000012A;
assign Y[4'b0100] [43] = 64'h00000000000004EA;
assign u[4'b0100] [43] = 64'h00000000000008EA;
assign v[4'b0100] [43] = 64'h0000000000000CEA;
assign X[4'b0100] [44] = 64'h000000000000012B;
assign Y[4'b0100] [44] = 64'h00000000000004EB;
assign u[4'b0100] [44] = 64'h00000000000008EB;
assign v[4'b0100] [44] = 64'h0000000000000CEB;
assign X[4'b0100] [45] = 64'h000000000000012C;
assign Y[4'b0100] [45] = 64'h00000000000004EC;
assign u[4'b0100] [45] = 64'h00000000000008EC;
assign v[4'b0100] [45] = 64'h0000000000000CEC;
assign X[4'b0100] [46] = 64'h000000000000012D;
assign Y[4'b0100] [46] = 64'h00000000000004ED;
assign u[4'b0100] [46] = 64'h00000000000008ED;
assign v[4'b0100] [46] = 64'h0000000000000CED;
assign X[4'b0100] [47] = 64'h000000000000012E;
assign Y[4'b0100] [47] = 64'h00000000000004EE;
assign u[4'b0100] [47] = 64'h00000000000008EE;
assign v[4'b0100] [47] = 64'h0000000000000CEE;
assign X[4'b0100] [48] = 64'h000000000000012F;
assign Y[4'b0100] [48] = 64'h00000000000004EF;
assign u[4'b0100] [48] = 64'h00000000000008EF;
assign v[4'b0100] [48] = 64'h0000000000000CEF;
assign X[4'b0100] [49] = 64'h0000000000000130;
assign Y[4'b0100] [49] = 64'h00000000000004F0;
assign u[4'b0100] [49] = 64'h00000000000008F0;
assign v[4'b0100] [49] = 64'h0000000000000CF0;
assign X[4'b0100] [50] = 64'h0000000000000131;
assign Y[4'b0100] [50] = 64'h00000000000004F1;
assign u[4'b0100] [50] = 64'h00000000000008F1;
assign v[4'b0100] [50] = 64'h0000000000000CF1;
assign X[4'b0100] [51] = 64'h0000000000000132;
assign Y[4'b0100] [51] = 64'h00000000000004F2;
assign u[4'b0100] [51] = 64'h00000000000008F2;
assign v[4'b0100] [51] = 64'h0000000000000CF2;
assign X[4'b0100] [52] = 64'h0000000000000133;
assign Y[4'b0100] [52] = 64'h00000000000004F3;
assign u[4'b0100] [52] = 64'h00000000000008F3;
assign v[4'b0100] [52] = 64'h0000000000000CF3;
assign X[4'b0100] [53] = 64'h0000000000000134;
assign Y[4'b0100] [53] = 64'h00000000000004F4;
assign u[4'b0100] [53] = 64'h00000000000008F4;
assign v[4'b0100] [53] = 64'h0000000000000CF4;
assign X[4'b0100] [54] = 64'h0000000000000135;
assign Y[4'b0100] [54] = 64'h00000000000004F5;
assign u[4'b0100] [54] = 64'h00000000000008F5;
assign v[4'b0100] [54] = 64'h0000000000000CF5;
assign X[4'b0100] [55] = 64'h0000000000000136;
assign Y[4'b0100] [55] = 64'h00000000000004F6;
assign u[4'b0100] [55] = 64'h00000000000008F6;
assign v[4'b0100] [55] = 64'h0000000000000CF6;
assign X[4'b0100] [56] = 64'h0000000000000137;
assign Y[4'b0100] [56] = 64'h00000000000004F7;
assign u[4'b0100] [56] = 64'h00000000000008F7;
assign v[4'b0100] [56] = 64'h0000000000000CF7;
assign X[4'b0100] [57] = 64'h0000000000000138;
assign Y[4'b0100] [57] = 64'h00000000000004F8;
assign u[4'b0100] [57] = 64'h00000000000008F8;
assign v[4'b0100] [57] = 64'h0000000000000CF8;
assign X[4'b0100] [58] = 64'h0000000000000139;
assign Y[4'b0100] [58] = 64'h00000000000004F9;
assign u[4'b0100] [58] = 64'h00000000000008F9;
assign v[4'b0100] [58] = 64'h0000000000000CF9;
assign X[4'b0100] [59] = 64'h000000000000013A;
assign Y[4'b0100] [59] = 64'h00000000000004FA;
assign u[4'b0100] [59] = 64'h00000000000008FA;
assign v[4'b0100] [59] = 64'h0000000000000CFA;
assign X[4'b0100] [60] = 64'h000000000000013B;
assign Y[4'b0100] [60] = 64'h00000000000004FB;
assign u[4'b0100] [60] = 64'h00000000000008FB;
assign v[4'b0100] [60] = 64'h0000000000000CFB;
assign X[4'b0100] [61] = 64'h000000000000013C;
assign Y[4'b0100] [61] = 64'h00000000000004FC;
assign u[4'b0100] [61] = 64'h00000000000008FC;
assign v[4'b0100] [61] = 64'h0000000000000CFC;
assign X[4'b0100] [62] = 64'h000000000000013D;
assign Y[4'b0100] [62] = 64'h00000000000004FD;
assign u[4'b0100] [62] = 64'h00000000000008FD;
assign v[4'b0100] [62] = 64'h0000000000000CFD;
assign X[4'b0100] [63] = 64'h000000000000013E;
assign Y[4'b0100] [63] = 64'h00000000000004FE;
assign u[4'b0100] [63] = 64'h00000000000008FE;
assign v[4'b0100] [63] = 64'h0000000000000CFE;
assign X[4'b0100] [64] = 64'h000000000000013F;
assign Y[4'b0100] [64] = 64'h00000000000004FF;
assign u[4'b0100] [64] = 64'h00000000000008FF;
assign v[4'b0100] [64] = 64'h0000000000000CFF;
assign X[4'b0101] [01] = 64'h0000000000000140;
assign Y[4'b0101] [01] = 64'h0000000000000500;
assign u[4'b0101] [01] = 64'h0000000000000900;
assign v[4'b0101] [01] = 64'h0000000000000D00;
assign X[4'b0101] [02] = 64'h0000000000000141;
assign Y[4'b0101] [02] = 64'h0000000000000501;
assign u[4'b0101] [02] = 64'h0000000000000901;
assign v[4'b0101] [02] = 64'h0000000000000D01;
assign X[4'b0101] [03] = 64'h0000000000000142;
assign Y[4'b0101] [03] = 64'h0000000000000502;
assign u[4'b0101] [03] = 64'h0000000000000902;
assign v[4'b0101] [03] = 64'h0000000000000D02;
assign X[4'b0101] [04] = 64'h0000000000000143;
assign Y[4'b0101] [04] = 64'h0000000000000503;
assign u[4'b0101] [04] = 64'h0000000000000903;
assign v[4'b0101] [04] = 64'h0000000000000D03;
assign X[4'b0101] [05] = 64'h0000000000000144;
assign Y[4'b0101] [05] = 64'h0000000000000504;
assign u[4'b0101] [05] = 64'h0000000000000904;
assign v[4'b0101] [05] = 64'h0000000000000D04;
assign X[4'b0101] [06] = 64'h0000000000000145;
assign Y[4'b0101] [06] = 64'h0000000000000505;
assign u[4'b0101] [06] = 64'h0000000000000905;
assign v[4'b0101] [06] = 64'h0000000000000D05;
assign X[4'b0101] [07] = 64'h0000000000000146;
assign Y[4'b0101] [07] = 64'h0000000000000506;
assign u[4'b0101] [07] = 64'h0000000000000906;
assign v[4'b0101] [07] = 64'h0000000000000D06;
assign X[4'b0101] [08] = 64'h0000000000000147;
assign Y[4'b0101] [08] = 64'h0000000000000507;
assign u[4'b0101] [08] = 64'h0000000000000907;
assign v[4'b0101] [08] = 64'h0000000000000D07;
assign X[4'b0101] [09] = 64'h0000000000000148;
assign Y[4'b0101] [09] = 64'h0000000000000508;
assign u[4'b0101] [09] = 64'h0000000000000908;
assign v[4'b0101] [09] = 64'h0000000000000D08;
assign X[4'b0101] [10] = 64'h0000000000000149;
assign Y[4'b0101] [10] = 64'h0000000000000509;
assign u[4'b0101] [10] = 64'h0000000000000909;
assign v[4'b0101] [10] = 64'h0000000000000D09;
assign X[4'b0101] [11] = 64'h000000000000014A;
assign Y[4'b0101] [11] = 64'h000000000000050A;
assign u[4'b0101] [11] = 64'h000000000000090A;
assign v[4'b0101] [11] = 64'h0000000000000D0A;
assign X[4'b0101] [12] = 64'h000000000000014B;
assign Y[4'b0101] [12] = 64'h000000000000050B;
assign u[4'b0101] [12] = 64'h000000000000090B;
assign v[4'b0101] [12] = 64'h0000000000000D0B;
assign X[4'b0101] [13] = 64'h000000000000014C;
assign Y[4'b0101] [13] = 64'h000000000000050C;
assign u[4'b0101] [13] = 64'h000000000000090C;
assign v[4'b0101] [13] = 64'h0000000000000D0C;
assign X[4'b0101] [14] = 64'h000000000000014D;
assign Y[4'b0101] [14] = 64'h000000000000050D;
assign u[4'b0101] [14] = 64'h000000000000090D;
assign v[4'b0101] [14] = 64'h0000000000000D0D;
assign X[4'b0101] [15] = 64'h000000000000014E;
assign Y[4'b0101] [15] = 64'h000000000000050E;
assign u[4'b0101] [15] = 64'h000000000000090E;
assign v[4'b0101] [15] = 64'h0000000000000D0E;
assign X[4'b0101] [16] = 64'h000000000000014F;
assign Y[4'b0101] [16] = 64'h000000000000050F;
assign u[4'b0101] [16] = 64'h000000000000090F;
assign v[4'b0101] [16] = 64'h0000000000000D0F;
assign X[4'b0101] [17] = 64'h0000000000000150;
assign Y[4'b0101] [17] = 64'h0000000000000510;
assign u[4'b0101] [17] = 64'h0000000000000910;
assign v[4'b0101] [17] = 64'h0000000000000D10;
assign X[4'b0101] [18] = 64'h0000000000000151;
assign Y[4'b0101] [18] = 64'h0000000000000511;
assign u[4'b0101] [18] = 64'h0000000000000911;
assign v[4'b0101] [18] = 64'h0000000000000D11;
assign X[4'b0101] [19] = 64'h0000000000000152;
assign Y[4'b0101] [19] = 64'h0000000000000512;
assign u[4'b0101] [19] = 64'h0000000000000912;
assign v[4'b0101] [19] = 64'h0000000000000D12;
assign X[4'b0101] [20] = 64'h0000000000000153;
assign Y[4'b0101] [20] = 64'h0000000000000513;
assign u[4'b0101] [20] = 64'h0000000000000913;
assign v[4'b0101] [20] = 64'h0000000000000D13;
assign X[4'b0101] [21] = 64'h0000000000000154;
assign Y[4'b0101] [21] = 64'h0000000000000514;
assign u[4'b0101] [21] = 64'h0000000000000914;
assign v[4'b0101] [21] = 64'h0000000000000D14;
assign X[4'b0101] [22] = 64'h0000000000000155;
assign Y[4'b0101] [22] = 64'h0000000000000515;
assign u[4'b0101] [22] = 64'h0000000000000915;
assign v[4'b0101] [22] = 64'h0000000000000D15;
assign X[4'b0101] [23] = 64'h0000000000000156;
assign Y[4'b0101] [23] = 64'h0000000000000516;
assign u[4'b0101] [23] = 64'h0000000000000916;
assign v[4'b0101] [23] = 64'h0000000000000D16;
assign X[4'b0101] [24] = 64'h0000000000000157;
assign Y[4'b0101] [24] = 64'h0000000000000517;
assign u[4'b0101] [24] = 64'h0000000000000917;
assign v[4'b0101] [24] = 64'h0000000000000D17;
assign X[4'b0101] [25] = 64'h0000000000000158;
assign Y[4'b0101] [25] = 64'h0000000000000518;
assign u[4'b0101] [25] = 64'h0000000000000918;
assign v[4'b0101] [25] = 64'h0000000000000D18;
assign X[4'b0101] [26] = 64'h0000000000000159;
assign Y[4'b0101] [26] = 64'h0000000000000519;
assign u[4'b0101] [26] = 64'h0000000000000919;
assign v[4'b0101] [26] = 64'h0000000000000D19;
assign X[4'b0101] [27] = 64'h000000000000015A;
assign Y[4'b0101] [27] = 64'h000000000000051A;
assign u[4'b0101] [27] = 64'h000000000000091A;
assign v[4'b0101] [27] = 64'h0000000000000D1A;
assign X[4'b0101] [28] = 64'h000000000000015B;
assign Y[4'b0101] [28] = 64'h000000000000051B;
assign u[4'b0101] [28] = 64'h000000000000091B;
assign v[4'b0101] [28] = 64'h0000000000000D1B;
assign X[4'b0101] [29] = 64'h000000000000015C;
assign Y[4'b0101] [29] = 64'h000000000000051C;
assign u[4'b0101] [29] = 64'h000000000000091C;
assign v[4'b0101] [29] = 64'h0000000000000D1C;
assign X[4'b0101] [30] = 64'h000000000000015D;
assign Y[4'b0101] [30] = 64'h000000000000051D;
assign u[4'b0101] [30] = 64'h000000000000091D;
assign v[4'b0101] [30] = 64'h0000000000000D1D;
assign X[4'b0101] [31] = 64'h000000000000015E;
assign Y[4'b0101] [31] = 64'h000000000000051E;
assign u[4'b0101] [31] = 64'h000000000000091E;
assign v[4'b0101] [31] = 64'h0000000000000D1E;
assign X[4'b0101] [32] = 64'h000000000000015F;
assign Y[4'b0101] [32] = 64'h000000000000051F;
assign u[4'b0101] [32] = 64'h000000000000091F;
assign v[4'b0101] [32] = 64'h0000000000000D1F;
assign X[4'b0101] [33] = 64'h0000000000000160;
assign Y[4'b0101] [33] = 64'h0000000000000520;
assign u[4'b0101] [33] = 64'h0000000000000920;
assign v[4'b0101] [33] = 64'h0000000000000D20;
assign X[4'b0101] [34] = 64'h0000000000000161;
assign Y[4'b0101] [34] = 64'h0000000000000521;
assign u[4'b0101] [34] = 64'h0000000000000921;
assign v[4'b0101] [34] = 64'h0000000000000D21;
assign X[4'b0101] [35] = 64'h0000000000000162;
assign Y[4'b0101] [35] = 64'h0000000000000522;
assign u[4'b0101] [35] = 64'h0000000000000922;
assign v[4'b0101] [35] = 64'h0000000000000D22;
assign X[4'b0101] [36] = 64'h0000000000000163;
assign Y[4'b0101] [36] = 64'h0000000000000523;
assign u[4'b0101] [36] = 64'h0000000000000923;
assign v[4'b0101] [36] = 64'h0000000000000D23;
assign X[4'b0101] [37] = 64'h0000000000000164;
assign Y[4'b0101] [37] = 64'h0000000000000524;
assign u[4'b0101] [37] = 64'h0000000000000924;
assign v[4'b0101] [37] = 64'h0000000000000D24;
assign X[4'b0101] [38] = 64'h0000000000000165;
assign Y[4'b0101] [38] = 64'h0000000000000525;
assign u[4'b0101] [38] = 64'h0000000000000925;
assign v[4'b0101] [38] = 64'h0000000000000D25;
assign X[4'b0101] [39] = 64'h0000000000000166;
assign Y[4'b0101] [39] = 64'h0000000000000526;
assign u[4'b0101] [39] = 64'h0000000000000926;
assign v[4'b0101] [39] = 64'h0000000000000D26;
assign X[4'b0101] [40] = 64'h0000000000000167;
assign Y[4'b0101] [40] = 64'h0000000000000527;
assign u[4'b0101] [40] = 64'h0000000000000927;
assign v[4'b0101] [40] = 64'h0000000000000D27;
assign X[4'b0101] [41] = 64'h0000000000000168;
assign Y[4'b0101] [41] = 64'h0000000000000528;
assign u[4'b0101] [41] = 64'h0000000000000928;
assign v[4'b0101] [41] = 64'h0000000000000D28;
assign X[4'b0101] [42] = 64'h0000000000000169;
assign Y[4'b0101] [42] = 64'h0000000000000529;
assign u[4'b0101] [42] = 64'h0000000000000929;
assign v[4'b0101] [42] = 64'h0000000000000D29;
assign X[4'b0101] [43] = 64'h000000000000016A;
assign Y[4'b0101] [43] = 64'h000000000000052A;
assign u[4'b0101] [43] = 64'h000000000000092A;
assign v[4'b0101] [43] = 64'h0000000000000D2A;
assign X[4'b0101] [44] = 64'h000000000000016B;
assign Y[4'b0101] [44] = 64'h000000000000052B;
assign u[4'b0101] [44] = 64'h000000000000092B;
assign v[4'b0101] [44] = 64'h0000000000000D2B;
assign X[4'b0101] [45] = 64'h000000000000016C;
assign Y[4'b0101] [45] = 64'h000000000000052C;
assign u[4'b0101] [45] = 64'h000000000000092C;
assign v[4'b0101] [45] = 64'h0000000000000D2C;
assign X[4'b0101] [46] = 64'h000000000000016D;
assign Y[4'b0101] [46] = 64'h000000000000052D;
assign u[4'b0101] [46] = 64'h000000000000092D;
assign v[4'b0101] [46] = 64'h0000000000000D2D;
assign X[4'b0101] [47] = 64'h000000000000016E;
assign Y[4'b0101] [47] = 64'h000000000000052E;
assign u[4'b0101] [47] = 64'h000000000000092E;
assign v[4'b0101] [47] = 64'h0000000000000D2E;
assign X[4'b0101] [48] = 64'h000000000000016F;
assign Y[4'b0101] [48] = 64'h000000000000052F;
assign u[4'b0101] [48] = 64'h000000000000092F;
assign v[4'b0101] [48] = 64'h0000000000000D2F;
assign X[4'b0101] [49] = 64'h0000000000000170;
assign Y[4'b0101] [49] = 64'h0000000000000530;
assign u[4'b0101] [49] = 64'h0000000000000930;
assign v[4'b0101] [49] = 64'h0000000000000D30;
assign X[4'b0101] [50] = 64'h0000000000000171;
assign Y[4'b0101] [50] = 64'h0000000000000531;
assign u[4'b0101] [50] = 64'h0000000000000931;
assign v[4'b0101] [50] = 64'h0000000000000D31;
assign X[4'b0101] [51] = 64'h0000000000000172;
assign Y[4'b0101] [51] = 64'h0000000000000532;
assign u[4'b0101] [51] = 64'h0000000000000932;
assign v[4'b0101] [51] = 64'h0000000000000D32;
assign X[4'b0101] [52] = 64'h0000000000000173;
assign Y[4'b0101] [52] = 64'h0000000000000533;
assign u[4'b0101] [52] = 64'h0000000000000933;
assign v[4'b0101] [52] = 64'h0000000000000D33;
assign X[4'b0101] [53] = 64'h0000000000000174;
assign Y[4'b0101] [53] = 64'h0000000000000534;
assign u[4'b0101] [53] = 64'h0000000000000934;
assign v[4'b0101] [53] = 64'h0000000000000D34;
assign X[4'b0101] [54] = 64'h0000000000000175;
assign Y[4'b0101] [54] = 64'h0000000000000535;
assign u[4'b0101] [54] = 64'h0000000000000935;
assign v[4'b0101] [54] = 64'h0000000000000D35;
assign X[4'b0101] [55] = 64'h0000000000000176;
assign Y[4'b0101] [55] = 64'h0000000000000536;
assign u[4'b0101] [55] = 64'h0000000000000936;
assign v[4'b0101] [55] = 64'h0000000000000D36;
assign X[4'b0101] [56] = 64'h0000000000000177;
assign Y[4'b0101] [56] = 64'h0000000000000537;
assign u[4'b0101] [56] = 64'h0000000000000937;
assign v[4'b0101] [56] = 64'h0000000000000D37;
assign X[4'b0101] [57] = 64'h0000000000000178;
assign Y[4'b0101] [57] = 64'h0000000000000538;
assign u[4'b0101] [57] = 64'h0000000000000938;
assign v[4'b0101] [57] = 64'h0000000000000D38;
assign X[4'b0101] [58] = 64'h0000000000000179;
assign Y[4'b0101] [58] = 64'h0000000000000539;
assign u[4'b0101] [58] = 64'h0000000000000939;
assign v[4'b0101] [58] = 64'h0000000000000D39;
assign X[4'b0101] [59] = 64'h000000000000017A;
assign Y[4'b0101] [59] = 64'h000000000000053A;
assign u[4'b0101] [59] = 64'h000000000000093A;
assign v[4'b0101] [59] = 64'h0000000000000D3A;
assign X[4'b0101] [60] = 64'h000000000000017B;
assign Y[4'b0101] [60] = 64'h000000000000053B;
assign u[4'b0101] [60] = 64'h000000000000093B;
assign v[4'b0101] [60] = 64'h0000000000000D3B;
assign X[4'b0101] [61] = 64'h000000000000017C;
assign Y[4'b0101] [61] = 64'h000000000000053C;
assign u[4'b0101] [61] = 64'h000000000000093C;
assign v[4'b0101] [61] = 64'h0000000000000D3C;
assign X[4'b0101] [62] = 64'h000000000000017D;
assign Y[4'b0101] [62] = 64'h000000000000053D;
assign u[4'b0101] [62] = 64'h000000000000093D;
assign v[4'b0101] [62] = 64'h0000000000000D3D;
assign X[4'b0101] [63] = 64'h000000000000017E;
assign Y[4'b0101] [63] = 64'h000000000000053E;
assign u[4'b0101] [63] = 64'h000000000000093E;
assign v[4'b0101] [63] = 64'h0000000000000D3E;
assign X[4'b0101] [64] = 64'h000000000000017F;
assign Y[4'b0101] [64] = 64'h000000000000053F;
assign u[4'b0101] [64] = 64'h000000000000093F;
assign v[4'b0101] [64] = 64'h0000000000000D3F;
assign X[4'b0110] [01] = 64'h0000000000000180;
assign Y[4'b0110] [01] = 64'h0000000000000540;
assign u[4'b0110] [01] = 64'h0000000000000940;
assign v[4'b0110] [01] = 64'h0000000000000D40;
assign X[4'b0110] [02] = 64'h0000000000000181;
assign Y[4'b0110] [02] = 64'h0000000000000541;
assign u[4'b0110] [02] = 64'h0000000000000941;
assign v[4'b0110] [02] = 64'h0000000000000D41;
assign X[4'b0110] [03] = 64'h0000000000000182;
assign Y[4'b0110] [03] = 64'h0000000000000542;
assign u[4'b0110] [03] = 64'h0000000000000942;
assign v[4'b0110] [03] = 64'h0000000000000D42;
assign X[4'b0110] [04] = 64'h0000000000000183;
assign Y[4'b0110] [04] = 64'h0000000000000543;
assign u[4'b0110] [04] = 64'h0000000000000943;
assign v[4'b0110] [04] = 64'h0000000000000D43;
assign X[4'b0110] [05] = 64'h0000000000000184;
assign Y[4'b0110] [05] = 64'h0000000000000544;
assign u[4'b0110] [05] = 64'h0000000000000944;
assign v[4'b0110] [05] = 64'h0000000000000D44;
assign X[4'b0110] [06] = 64'h0000000000000185;
assign Y[4'b0110] [06] = 64'h0000000000000545;
assign u[4'b0110] [06] = 64'h0000000000000945;
assign v[4'b0110] [06] = 64'h0000000000000D45;
assign X[4'b0110] [07] = 64'h0000000000000186;
assign Y[4'b0110] [07] = 64'h0000000000000546;
assign u[4'b0110] [07] = 64'h0000000000000946;
assign v[4'b0110] [07] = 64'h0000000000000D46;
assign X[4'b0110] [08] = 64'h0000000000000187;
assign Y[4'b0110] [08] = 64'h0000000000000547;
assign u[4'b0110] [08] = 64'h0000000000000947;
assign v[4'b0110] [08] = 64'h0000000000000D47;
assign X[4'b0110] [09] = 64'h0000000000000188;
assign Y[4'b0110] [09] = 64'h0000000000000548;
assign u[4'b0110] [09] = 64'h0000000000000948;
assign v[4'b0110] [09] = 64'h0000000000000D48;
assign X[4'b0110] [10] = 64'h0000000000000189;
assign Y[4'b0110] [10] = 64'h0000000000000549;
assign u[4'b0110] [10] = 64'h0000000000000949;
assign v[4'b0110] [10] = 64'h0000000000000D49;
assign X[4'b0110] [11] = 64'h000000000000018A;
assign Y[4'b0110] [11] = 64'h000000000000054A;
assign u[4'b0110] [11] = 64'h000000000000094A;
assign v[4'b0110] [11] = 64'h0000000000000D4A;
assign X[4'b0110] [12] = 64'h000000000000018B;
assign Y[4'b0110] [12] = 64'h000000000000054B;
assign u[4'b0110] [12] = 64'h000000000000094B;
assign v[4'b0110] [12] = 64'h0000000000000D4B;
assign X[4'b0110] [13] = 64'h000000000000018C;
assign Y[4'b0110] [13] = 64'h000000000000054C;
assign u[4'b0110] [13] = 64'h000000000000094C;
assign v[4'b0110] [13] = 64'h0000000000000D4C;
assign X[4'b0110] [14] = 64'h000000000000018D;
assign Y[4'b0110] [14] = 64'h000000000000054D;
assign u[4'b0110] [14] = 64'h000000000000094D;
assign v[4'b0110] [14] = 64'h0000000000000D4D;
assign X[4'b0110] [15] = 64'h000000000000018E;
assign Y[4'b0110] [15] = 64'h000000000000054E;
assign u[4'b0110] [15] = 64'h000000000000094E;
assign v[4'b0110] [15] = 64'h0000000000000D4E;
assign X[4'b0110] [16] = 64'h000000000000018F;
assign Y[4'b0110] [16] = 64'h000000000000054F;
assign u[4'b0110] [16] = 64'h000000000000094F;
assign v[4'b0110] [16] = 64'h0000000000000D4F;
assign X[4'b0110] [17] = 64'h0000000000000190;
assign Y[4'b0110] [17] = 64'h0000000000000550;
assign u[4'b0110] [17] = 64'h0000000000000950;
assign v[4'b0110] [17] = 64'h0000000000000D50;
assign X[4'b0110] [18] = 64'h0000000000000191;
assign Y[4'b0110] [18] = 64'h0000000000000551;
assign u[4'b0110] [18] = 64'h0000000000000951;
assign v[4'b0110] [18] = 64'h0000000000000D51;
assign X[4'b0110] [19] = 64'h0000000000000192;
assign Y[4'b0110] [19] = 64'h0000000000000552;
assign u[4'b0110] [19] = 64'h0000000000000952;
assign v[4'b0110] [19] = 64'h0000000000000D52;
assign X[4'b0110] [20] = 64'h0000000000000193;
assign Y[4'b0110] [20] = 64'h0000000000000553;
assign u[4'b0110] [20] = 64'h0000000000000953;
assign v[4'b0110] [20] = 64'h0000000000000D53;
assign X[4'b0110] [21] = 64'h0000000000000194;
assign Y[4'b0110] [21] = 64'h0000000000000554;
assign u[4'b0110] [21] = 64'h0000000000000954;
assign v[4'b0110] [21] = 64'h0000000000000D54;
assign X[4'b0110] [22] = 64'h0000000000000195;
assign Y[4'b0110] [22] = 64'h0000000000000555;
assign u[4'b0110] [22] = 64'h0000000000000955;
assign v[4'b0110] [22] = 64'h0000000000000D55;
assign X[4'b0110] [23] = 64'h0000000000000196;
assign Y[4'b0110] [23] = 64'h0000000000000556;
assign u[4'b0110] [23] = 64'h0000000000000956;
assign v[4'b0110] [23] = 64'h0000000000000D56;
assign X[4'b0110] [24] = 64'h0000000000000197;
assign Y[4'b0110] [24] = 64'h0000000000000557;
assign u[4'b0110] [24] = 64'h0000000000000957;
assign v[4'b0110] [24] = 64'h0000000000000D57;
assign X[4'b0110] [25] = 64'h0000000000000198;
assign Y[4'b0110] [25] = 64'h0000000000000558;
assign u[4'b0110] [25] = 64'h0000000000000958;
assign v[4'b0110] [25] = 64'h0000000000000D58;
assign X[4'b0110] [26] = 64'h0000000000000199;
assign Y[4'b0110] [26] = 64'h0000000000000559;
assign u[4'b0110] [26] = 64'h0000000000000959;
assign v[4'b0110] [26] = 64'h0000000000000D59;
assign X[4'b0110] [27] = 64'h000000000000019A;
assign Y[4'b0110] [27] = 64'h000000000000055A;
assign u[4'b0110] [27] = 64'h000000000000095A;
assign v[4'b0110] [27] = 64'h0000000000000D5A;
assign X[4'b0110] [28] = 64'h000000000000019B;
assign Y[4'b0110] [28] = 64'h000000000000055B;
assign u[4'b0110] [28] = 64'h000000000000095B;
assign v[4'b0110] [28] = 64'h0000000000000D5B;
assign X[4'b0110] [29] = 64'h000000000000019C;
assign Y[4'b0110] [29] = 64'h000000000000055C;
assign u[4'b0110] [29] = 64'h000000000000095C;
assign v[4'b0110] [29] = 64'h0000000000000D5C;
assign X[4'b0110] [30] = 64'h000000000000019D;
assign Y[4'b0110] [30] = 64'h000000000000055D;
assign u[4'b0110] [30] = 64'h000000000000095D;
assign v[4'b0110] [30] = 64'h0000000000000D5D;
assign X[4'b0110] [31] = 64'h000000000000019E;
assign Y[4'b0110] [31] = 64'h000000000000055E;
assign u[4'b0110] [31] = 64'h000000000000095E;
assign v[4'b0110] [31] = 64'h0000000000000D5E;
assign X[4'b0110] [32] = 64'h000000000000019F;
assign Y[4'b0110] [32] = 64'h000000000000055F;
assign u[4'b0110] [32] = 64'h000000000000095F;
assign v[4'b0110] [32] = 64'h0000000000000D5F;
assign X[4'b0110] [33] = 64'h00000000000001A0;
assign Y[4'b0110] [33] = 64'h0000000000000560;
assign u[4'b0110] [33] = 64'h0000000000000960;
assign v[4'b0110] [33] = 64'h0000000000000D60;
assign X[4'b0110] [34] = 64'h00000000000001A1;
assign Y[4'b0110] [34] = 64'h0000000000000561;
assign u[4'b0110] [34] = 64'h0000000000000961;
assign v[4'b0110] [34] = 64'h0000000000000D61;
assign X[4'b0110] [35] = 64'h00000000000001A2;
assign Y[4'b0110] [35] = 64'h0000000000000562;
assign u[4'b0110] [35] = 64'h0000000000000962;
assign v[4'b0110] [35] = 64'h0000000000000D62;
assign X[4'b0110] [36] = 64'h00000000000001A3;
assign Y[4'b0110] [36] = 64'h0000000000000563;
assign u[4'b0110] [36] = 64'h0000000000000963;
assign v[4'b0110] [36] = 64'h0000000000000D63;
assign X[4'b0110] [37] = 64'h00000000000001A4;
assign Y[4'b0110] [37] = 64'h0000000000000564;
assign u[4'b0110] [37] = 64'h0000000000000964;
assign v[4'b0110] [37] = 64'h0000000000000D64;
assign X[4'b0110] [38] = 64'h00000000000001A5;
assign Y[4'b0110] [38] = 64'h0000000000000565;
assign u[4'b0110] [38] = 64'h0000000000000965;
assign v[4'b0110] [38] = 64'h0000000000000D65;
assign X[4'b0110] [39] = 64'h00000000000001A6;
assign Y[4'b0110] [39] = 64'h0000000000000566;
assign u[4'b0110] [39] = 64'h0000000000000966;
assign v[4'b0110] [39] = 64'h0000000000000D66;
assign X[4'b0110] [40] = 64'h00000000000001A7;
assign Y[4'b0110] [40] = 64'h0000000000000567;
assign u[4'b0110] [40] = 64'h0000000000000967;
assign v[4'b0110] [40] = 64'h0000000000000D67;
assign X[4'b0110] [41] = 64'h00000000000001A8;
assign Y[4'b0110] [41] = 64'h0000000000000568;
assign u[4'b0110] [41] = 64'h0000000000000968;
assign v[4'b0110] [41] = 64'h0000000000000D68;
assign X[4'b0110] [42] = 64'h00000000000001A9;
assign Y[4'b0110] [42] = 64'h0000000000000569;
assign u[4'b0110] [42] = 64'h0000000000000969;
assign v[4'b0110] [42] = 64'h0000000000000D69;
assign X[4'b0110] [43] = 64'h00000000000001AA;
assign Y[4'b0110] [43] = 64'h000000000000056A;
assign u[4'b0110] [43] = 64'h000000000000096A;
assign v[4'b0110] [43] = 64'h0000000000000D6A;
assign X[4'b0110] [44] = 64'h00000000000001AB;
assign Y[4'b0110] [44] = 64'h000000000000056B;
assign u[4'b0110] [44] = 64'h000000000000096B;
assign v[4'b0110] [44] = 64'h0000000000000D6B;
assign X[4'b0110] [45] = 64'h00000000000001AC;
assign Y[4'b0110] [45] = 64'h000000000000056C;
assign u[4'b0110] [45] = 64'h000000000000096C;
assign v[4'b0110] [45] = 64'h0000000000000D6C;
assign X[4'b0110] [46] = 64'h00000000000001AD;
assign Y[4'b0110] [46] = 64'h000000000000056D;
assign u[4'b0110] [46] = 64'h000000000000096D;
assign v[4'b0110] [46] = 64'h0000000000000D6D;
assign X[4'b0110] [47] = 64'h00000000000001AE;
assign Y[4'b0110] [47] = 64'h000000000000056E;
assign u[4'b0110] [47] = 64'h000000000000096E;
assign v[4'b0110] [47] = 64'h0000000000000D6E;
assign X[4'b0110] [48] = 64'h00000000000001AF;
assign Y[4'b0110] [48] = 64'h000000000000056F;
assign u[4'b0110] [48] = 64'h000000000000096F;
assign v[4'b0110] [48] = 64'h0000000000000D6F;
assign X[4'b0110] [49] = 64'h00000000000001B0;
assign Y[4'b0110] [49] = 64'h0000000000000570;
assign u[4'b0110] [49] = 64'h0000000000000970;
assign v[4'b0110] [49] = 64'h0000000000000D70;
assign X[4'b0110] [50] = 64'h00000000000001B1;
assign Y[4'b0110] [50] = 64'h0000000000000571;
assign u[4'b0110] [50] = 64'h0000000000000971;
assign v[4'b0110] [50] = 64'h0000000000000D71;
assign X[4'b0110] [51] = 64'h00000000000001B2;
assign Y[4'b0110] [51] = 64'h0000000000000572;
assign u[4'b0110] [51] = 64'h0000000000000972;
assign v[4'b0110] [51] = 64'h0000000000000D72;
assign X[4'b0110] [52] = 64'h00000000000001B3;
assign Y[4'b0110] [52] = 64'h0000000000000573;
assign u[4'b0110] [52] = 64'h0000000000000973;
assign v[4'b0110] [52] = 64'h0000000000000D73;
assign X[4'b0110] [53] = 64'h00000000000001B4;
assign Y[4'b0110] [53] = 64'h0000000000000574;
assign u[4'b0110] [53] = 64'h0000000000000974;
assign v[4'b0110] [53] = 64'h0000000000000D74;
assign X[4'b0110] [54] = 64'h00000000000001B5;
assign Y[4'b0110] [54] = 64'h0000000000000575;
assign u[4'b0110] [54] = 64'h0000000000000975;
assign v[4'b0110] [54] = 64'h0000000000000D75;
assign X[4'b0110] [55] = 64'h00000000000001B6;
assign Y[4'b0110] [55] = 64'h0000000000000576;
assign u[4'b0110] [55] = 64'h0000000000000976;
assign v[4'b0110] [55] = 64'h0000000000000D76;
assign X[4'b0110] [56] = 64'h00000000000001B7;
assign Y[4'b0110] [56] = 64'h0000000000000577;
assign u[4'b0110] [56] = 64'h0000000000000977;
assign v[4'b0110] [56] = 64'h0000000000000D77;
assign X[4'b0110] [57] = 64'h00000000000001B8;
assign Y[4'b0110] [57] = 64'h0000000000000578;
assign u[4'b0110] [57] = 64'h0000000000000978;
assign v[4'b0110] [57] = 64'h0000000000000D78;
assign X[4'b0110] [58] = 64'h00000000000001B9;
assign Y[4'b0110] [58] = 64'h0000000000000579;
assign u[4'b0110] [58] = 64'h0000000000000979;
assign v[4'b0110] [58] = 64'h0000000000000D79;
assign X[4'b0110] [59] = 64'h00000000000001BA;
assign Y[4'b0110] [59] = 64'h000000000000057A;
assign u[4'b0110] [59] = 64'h000000000000097A;
assign v[4'b0110] [59] = 64'h0000000000000D7A;
assign X[4'b0110] [60] = 64'h00000000000001BB;
assign Y[4'b0110] [60] = 64'h000000000000057B;
assign u[4'b0110] [60] = 64'h000000000000097B;
assign v[4'b0110] [60] = 64'h0000000000000D7B;
assign X[4'b0110] [61] = 64'h00000000000001BC;
assign Y[4'b0110] [61] = 64'h000000000000057C;
assign u[4'b0110] [61] = 64'h000000000000097C;
assign v[4'b0110] [61] = 64'h0000000000000D7C;
assign X[4'b0110] [62] = 64'h00000000000001BD;
assign Y[4'b0110] [62] = 64'h000000000000057D;
assign u[4'b0110] [62] = 64'h000000000000097D;
assign v[4'b0110] [62] = 64'h0000000000000D7D;
assign X[4'b0110] [63] = 64'h00000000000001BE;
assign Y[4'b0110] [63] = 64'h000000000000057E;
assign u[4'b0110] [63] = 64'h000000000000097E;
assign v[4'b0110] [63] = 64'h0000000000000D7E;
assign X[4'b0110] [64] = 64'h00000000000001BF;
assign Y[4'b0110] [64] = 64'h000000000000057F;
assign u[4'b0110] [64] = 64'h000000000000097F;
assign v[4'b0110] [64] = 64'h0000000000000D7F;
assign X[4'b0111] [01] = 64'h00000000000001C0;
assign Y[4'b0111] [01] = 64'h0000000000000580;
assign u[4'b0111] [01] = 64'h0000000000000980;
assign v[4'b0111] [01] = 64'h0000000000000D80;
assign X[4'b0111] [02] = 64'h00000000000001C1;
assign Y[4'b0111] [02] = 64'h0000000000000581;
assign u[4'b0111] [02] = 64'h0000000000000981;
assign v[4'b0111] [02] = 64'h0000000000000D81;
assign X[4'b0111] [03] = 64'h00000000000001C2;
assign Y[4'b0111] [03] = 64'h0000000000000582;
assign u[4'b0111] [03] = 64'h0000000000000982;
assign v[4'b0111] [03] = 64'h0000000000000D82;
assign X[4'b0111] [04] = 64'h00000000000001C3;
assign Y[4'b0111] [04] = 64'h0000000000000583;
assign u[4'b0111] [04] = 64'h0000000000000983;
assign v[4'b0111] [04] = 64'h0000000000000D83;
assign X[4'b0111] [05] = 64'h00000000000001C4;
assign Y[4'b0111] [05] = 64'h0000000000000584;
assign u[4'b0111] [05] = 64'h0000000000000984;
assign v[4'b0111] [05] = 64'h0000000000000D84;
assign X[4'b0111] [06] = 64'h00000000000001C5;
assign Y[4'b0111] [06] = 64'h0000000000000585;
assign u[4'b0111] [06] = 64'h0000000000000985;
assign v[4'b0111] [06] = 64'h0000000000000D85;
assign X[4'b0111] [07] = 64'h00000000000001C6;
assign Y[4'b0111] [07] = 64'h0000000000000586;
assign u[4'b0111] [07] = 64'h0000000000000986;
assign v[4'b0111] [07] = 64'h0000000000000D86;
assign X[4'b0111] [08] = 64'h00000000000001C7;
assign Y[4'b0111] [08] = 64'h0000000000000587;
assign u[4'b0111] [08] = 64'h0000000000000987;
assign v[4'b0111] [08] = 64'h0000000000000D87;
assign X[4'b0111] [09] = 64'h00000000000001C8;
assign Y[4'b0111] [09] = 64'h0000000000000588;
assign u[4'b0111] [09] = 64'h0000000000000988;
assign v[4'b0111] [09] = 64'h0000000000000D88;
assign X[4'b0111] [10] = 64'h00000000000001C9;
assign Y[4'b0111] [10] = 64'h0000000000000589;
assign u[4'b0111] [10] = 64'h0000000000000989;
assign v[4'b0111] [10] = 64'h0000000000000D89;
assign X[4'b0111] [11] = 64'h00000000000001CA;
assign Y[4'b0111] [11] = 64'h000000000000058A;
assign u[4'b0111] [11] = 64'h000000000000098A;
assign v[4'b0111] [11] = 64'h0000000000000D8A;
assign X[4'b0111] [12] = 64'h00000000000001CB;
assign Y[4'b0111] [12] = 64'h000000000000058B;
assign u[4'b0111] [12] = 64'h000000000000098B;
assign v[4'b0111] [12] = 64'h0000000000000D8B;
assign X[4'b0111] [13] = 64'h00000000000001CC;
assign Y[4'b0111] [13] = 64'h000000000000058C;
assign u[4'b0111] [13] = 64'h000000000000098C;
assign v[4'b0111] [13] = 64'h0000000000000D8C;
assign X[4'b0111] [14] = 64'h00000000000001CD;
assign Y[4'b0111] [14] = 64'h000000000000058D;
assign u[4'b0111] [14] = 64'h000000000000098D;
assign v[4'b0111] [14] = 64'h0000000000000D8D;
assign X[4'b0111] [15] = 64'h00000000000001CE;
assign Y[4'b0111] [15] = 64'h000000000000058E;
assign u[4'b0111] [15] = 64'h000000000000098E;
assign v[4'b0111] [15] = 64'h0000000000000D8E;
assign X[4'b0111] [16] = 64'h00000000000001CF;
assign Y[4'b0111] [16] = 64'h000000000000058F;
assign u[4'b0111] [16] = 64'h000000000000098F;
assign v[4'b0111] [16] = 64'h0000000000000D8F;
assign X[4'b0111] [17] = 64'h00000000000001D0;
assign Y[4'b0111] [17] = 64'h0000000000000590;
assign u[4'b0111] [17] = 64'h0000000000000990;
assign v[4'b0111] [17] = 64'h0000000000000D90;
assign X[4'b0111] [18] = 64'h00000000000001D1;
assign Y[4'b0111] [18] = 64'h0000000000000591;
assign u[4'b0111] [18] = 64'h0000000000000991;
assign v[4'b0111] [18] = 64'h0000000000000D91;
assign X[4'b0111] [19] = 64'h00000000000001D2;
assign Y[4'b0111] [19] = 64'h0000000000000592;
assign u[4'b0111] [19] = 64'h0000000000000992;
assign v[4'b0111] [19] = 64'h0000000000000D92;
assign X[4'b0111] [20] = 64'h00000000000001D3;
assign Y[4'b0111] [20] = 64'h0000000000000593;
assign u[4'b0111] [20] = 64'h0000000000000993;
assign v[4'b0111] [20] = 64'h0000000000000D93;
assign X[4'b0111] [21] = 64'h00000000000001D4;
assign Y[4'b0111] [21] = 64'h0000000000000594;
assign u[4'b0111] [21] = 64'h0000000000000994;
assign v[4'b0111] [21] = 64'h0000000000000D94;
assign X[4'b0111] [22] = 64'h00000000000001D5;
assign Y[4'b0111] [22] = 64'h0000000000000595;
assign u[4'b0111] [22] = 64'h0000000000000995;
assign v[4'b0111] [22] = 64'h0000000000000D95;
assign X[4'b0111] [23] = 64'h00000000000001D6;
assign Y[4'b0111] [23] = 64'h0000000000000596;
assign u[4'b0111] [23] = 64'h0000000000000996;
assign v[4'b0111] [23] = 64'h0000000000000D96;
assign X[4'b0111] [24] = 64'h00000000000001D7;
assign Y[4'b0111] [24] = 64'h0000000000000597;
assign u[4'b0111] [24] = 64'h0000000000000997;
assign v[4'b0111] [24] = 64'h0000000000000D97;
assign X[4'b0111] [25] = 64'h00000000000001D8;
assign Y[4'b0111] [25] = 64'h0000000000000598;
assign u[4'b0111] [25] = 64'h0000000000000998;
assign v[4'b0111] [25] = 64'h0000000000000D98;
assign X[4'b0111] [26] = 64'h00000000000001D9;
assign Y[4'b0111] [26] = 64'h0000000000000599;
assign u[4'b0111] [26] = 64'h0000000000000999;
assign v[4'b0111] [26] = 64'h0000000000000D99;
assign X[4'b0111] [27] = 64'h00000000000001DA;
assign Y[4'b0111] [27] = 64'h000000000000059A;
assign u[4'b0111] [27] = 64'h000000000000099A;
assign v[4'b0111] [27] = 64'h0000000000000D9A;
assign X[4'b0111] [28] = 64'h00000000000001DB;
assign Y[4'b0111] [28] = 64'h000000000000059B;
assign u[4'b0111] [28] = 64'h000000000000099B;
assign v[4'b0111] [28] = 64'h0000000000000D9B;
assign X[4'b0111] [29] = 64'h00000000000001DC;
assign Y[4'b0111] [29] = 64'h000000000000059C;
assign u[4'b0111] [29] = 64'h000000000000099C;
assign v[4'b0111] [29] = 64'h0000000000000D9C;
assign X[4'b0111] [30] = 64'h00000000000001DD;
assign Y[4'b0111] [30] = 64'h000000000000059D;
assign u[4'b0111] [30] = 64'h000000000000099D;
assign v[4'b0111] [30] = 64'h0000000000000D9D;
assign X[4'b0111] [31] = 64'h00000000000001DE;
assign Y[4'b0111] [31] = 64'h000000000000059E;
assign u[4'b0111] [31] = 64'h000000000000099E;
assign v[4'b0111] [31] = 64'h0000000000000D9E;
assign X[4'b0111] [32] = 64'h00000000000001DF;
assign Y[4'b0111] [32] = 64'h000000000000059F;
assign u[4'b0111] [32] = 64'h000000000000099F;
assign v[4'b0111] [32] = 64'h0000000000000D9F;
assign X[4'b0111] [33] = 64'h00000000000001E0;
assign Y[4'b0111] [33] = 64'h00000000000005A0;
assign u[4'b0111] [33] = 64'h00000000000009A0;
assign v[4'b0111] [33] = 64'h0000000000000DA0;
assign X[4'b0111] [34] = 64'h00000000000001E1;
assign Y[4'b0111] [34] = 64'h00000000000005A1;
assign u[4'b0111] [34] = 64'h00000000000009A1;
assign v[4'b0111] [34] = 64'h0000000000000DA1;
assign X[4'b0111] [35] = 64'h00000000000001E2;
assign Y[4'b0111] [35] = 64'h00000000000005A2;
assign u[4'b0111] [35] = 64'h00000000000009A2;
assign v[4'b0111] [35] = 64'h0000000000000DA2;
assign X[4'b0111] [36] = 64'h00000000000001E3;
assign Y[4'b0111] [36] = 64'h00000000000005A3;
assign u[4'b0111] [36] = 64'h00000000000009A3;
assign v[4'b0111] [36] = 64'h0000000000000DA3;
assign X[4'b0111] [37] = 64'h00000000000001E4;
assign Y[4'b0111] [37] = 64'h00000000000005A4;
assign u[4'b0111] [37] = 64'h00000000000009A4;
assign v[4'b0111] [37] = 64'h0000000000000DA4;
assign X[4'b0111] [38] = 64'h00000000000001E5;
assign Y[4'b0111] [38] = 64'h00000000000005A5;
assign u[4'b0111] [38] = 64'h00000000000009A5;
assign v[4'b0111] [38] = 64'h0000000000000DA5;
assign X[4'b0111] [39] = 64'h00000000000001E6;
assign Y[4'b0111] [39] = 64'h00000000000005A6;
assign u[4'b0111] [39] = 64'h00000000000009A6;
assign v[4'b0111] [39] = 64'h0000000000000DA6;
assign X[4'b0111] [40] = 64'h00000000000001E7;
assign Y[4'b0111] [40] = 64'h00000000000005A7;
assign u[4'b0111] [40] = 64'h00000000000009A7;
assign v[4'b0111] [40] = 64'h0000000000000DA7;
assign X[4'b0111] [41] = 64'h00000000000001E8;
assign Y[4'b0111] [41] = 64'h00000000000005A8;
assign u[4'b0111] [41] = 64'h00000000000009A8;
assign v[4'b0111] [41] = 64'h0000000000000DA8;
assign X[4'b0111] [42] = 64'h00000000000001E9;
assign Y[4'b0111] [42] = 64'h00000000000005A9;
assign u[4'b0111] [42] = 64'h00000000000009A9;
assign v[4'b0111] [42] = 64'h0000000000000DA9;
assign X[4'b0111] [43] = 64'h00000000000001EA;
assign Y[4'b0111] [43] = 64'h00000000000005AA;
assign u[4'b0111] [43] = 64'h00000000000009AA;
assign v[4'b0111] [43] = 64'h0000000000000DAA;
assign X[4'b0111] [44] = 64'h00000000000001EB;
assign Y[4'b0111] [44] = 64'h00000000000005AB;
assign u[4'b0111] [44] = 64'h00000000000009AB;
assign v[4'b0111] [44] = 64'h0000000000000DAB;
assign X[4'b0111] [45] = 64'h00000000000001EC;
assign Y[4'b0111] [45] = 64'h00000000000005AC;
assign u[4'b0111] [45] = 64'h00000000000009AC;
assign v[4'b0111] [45] = 64'h0000000000000DAC;
assign X[4'b0111] [46] = 64'h00000000000001ED;
assign Y[4'b0111] [46] = 64'h00000000000005AD;
assign u[4'b0111] [46] = 64'h00000000000009AD;
assign v[4'b0111] [46] = 64'h0000000000000DAD;
assign X[4'b0111] [47] = 64'h00000000000001EE;
assign Y[4'b0111] [47] = 64'h00000000000005AE;
assign u[4'b0111] [47] = 64'h00000000000009AE;
assign v[4'b0111] [47] = 64'h0000000000000DAE;
assign X[4'b0111] [48] = 64'h00000000000001EF;
assign Y[4'b0111] [48] = 64'h00000000000005AF;
assign u[4'b0111] [48] = 64'h00000000000009AF;
assign v[4'b0111] [48] = 64'h0000000000000DAF;
assign X[4'b0111] [49] = 64'h00000000000001F0;
assign Y[4'b0111] [49] = 64'h00000000000005B0;
assign u[4'b0111] [49] = 64'h00000000000009B0;
assign v[4'b0111] [49] = 64'h0000000000000DB0;
assign X[4'b0111] [50] = 64'h00000000000001F1;
assign Y[4'b0111] [50] = 64'h00000000000005B1;
assign u[4'b0111] [50] = 64'h00000000000009B1;
assign v[4'b0111] [50] = 64'h0000000000000DB1;
assign X[4'b0111] [51] = 64'h00000000000001F2;
assign Y[4'b0111] [51] = 64'h00000000000005B2;
assign u[4'b0111] [51] = 64'h00000000000009B2;
assign v[4'b0111] [51] = 64'h0000000000000DB2;
assign X[4'b0111] [52] = 64'h00000000000001F3;
assign Y[4'b0111] [52] = 64'h00000000000005B3;
assign u[4'b0111] [52] = 64'h00000000000009B3;
assign v[4'b0111] [52] = 64'h0000000000000DB3;
assign X[4'b0111] [53] = 64'h00000000000001F4;
assign Y[4'b0111] [53] = 64'h00000000000005B4;
assign u[4'b0111] [53] = 64'h00000000000009B4;
assign v[4'b0111] [53] = 64'h0000000000000DB4;
assign X[4'b0111] [54] = 64'h00000000000001F5;
assign Y[4'b0111] [54] = 64'h00000000000005B5;
assign u[4'b0111] [54] = 64'h00000000000009B5;
assign v[4'b0111] [54] = 64'h0000000000000DB5;
assign X[4'b0111] [55] = 64'h00000000000001F6;
assign Y[4'b0111] [55] = 64'h00000000000005B6;
assign u[4'b0111] [55] = 64'h00000000000009B6;
assign v[4'b0111] [55] = 64'h0000000000000DB6;
assign X[4'b0111] [56] = 64'h00000000000001F7;
assign Y[4'b0111] [56] = 64'h00000000000005B7;
assign u[4'b0111] [56] = 64'h00000000000009B7;
assign v[4'b0111] [56] = 64'h0000000000000DB7;
assign X[4'b0111] [57] = 64'h00000000000001F8;
assign Y[4'b0111] [57] = 64'h00000000000005B8;
assign u[4'b0111] [57] = 64'h00000000000009B8;
assign v[4'b0111] [57] = 64'h0000000000000DB8;
assign X[4'b0111] [58] = 64'h00000000000001F9;
assign Y[4'b0111] [58] = 64'h00000000000005B9;
assign u[4'b0111] [58] = 64'h00000000000009B9;
assign v[4'b0111] [58] = 64'h0000000000000DB9;
assign X[4'b0111] [59] = 64'h00000000000001FA;
assign Y[4'b0111] [59] = 64'h00000000000005BA;
assign u[4'b0111] [59] = 64'h00000000000009BA;
assign v[4'b0111] [59] = 64'h0000000000000DBA;
assign X[4'b0111] [60] = 64'h00000000000001FB;
assign Y[4'b0111] [60] = 64'h00000000000005BB;
assign u[4'b0111] [60] = 64'h00000000000009BB;
assign v[4'b0111] [60] = 64'h0000000000000DBB;
assign X[4'b0111] [61] = 64'h00000000000001FC;
assign Y[4'b0111] [61] = 64'h00000000000005BC;
assign u[4'b0111] [61] = 64'h00000000000009BC;
assign v[4'b0111] [61] = 64'h0000000000000DBC;
assign X[4'b0111] [62] = 64'h00000000000001FD;
assign Y[4'b0111] [62] = 64'h00000000000005BD;
assign u[4'b0111] [62] = 64'h00000000000009BD;
assign v[4'b0111] [62] = 64'h0000000000000DBD;
assign X[4'b0111] [63] = 64'h00000000000001FE;
assign Y[4'b0111] [63] = 64'h00000000000005BE;
assign u[4'b0111] [63] = 64'h00000000000009BE;
assign v[4'b0111] [63] = 64'h0000000000000DBE;
assign X[4'b0111] [64] = 64'h00000000000001FF;
assign Y[4'b0111] [64] = 64'h00000000000005BF;
assign u[4'b0111] [64] = 64'h00000000000009BF;
assign v[4'b0111] [64] = 64'h0000000000000DBF;
assign X[4'b1000] [01] = 64'h0000000000000200;
assign Y[4'b1000] [01] = 64'h00000000000005C0;
assign u[4'b1000] [01] = 64'h00000000000009C0;
assign v[4'b1000] [01] = 64'h0000000000000DC0;
assign X[4'b1000] [02] = 64'h0000000000000201;
assign Y[4'b1000] [02] = 64'h00000000000005C1;
assign u[4'b1000] [02] = 64'h00000000000009C1;
assign v[4'b1000] [02] = 64'h0000000000000DC1;
assign X[4'b1000] [03] = 64'h0000000000000202;
assign Y[4'b1000] [03] = 64'h00000000000005C2;
assign u[4'b1000] [03] = 64'h00000000000009C2;
assign v[4'b1000] [03] = 64'h0000000000000DC2;
assign X[4'b1000] [04] = 64'h0000000000000203;
assign Y[4'b1000] [04] = 64'h00000000000005C3;
assign u[4'b1000] [04] = 64'h00000000000009C3;
assign v[4'b1000] [04] = 64'h0000000000000DC3;
assign X[4'b1000] [05] = 64'h0000000000000204;
assign Y[4'b1000] [05] = 64'h00000000000005C4;
assign u[4'b1000] [05] = 64'h00000000000009C4;
assign v[4'b1000] [05] = 64'h0000000000000DC4;
assign X[4'b1000] [06] = 64'h0000000000000205;
assign Y[4'b1000] [06] = 64'h00000000000005C5;
assign u[4'b1000] [06] = 64'h00000000000009C5;
assign v[4'b1000] [06] = 64'h0000000000000DC5;
assign X[4'b1000] [07] = 64'h0000000000000206;
assign Y[4'b1000] [07] = 64'h00000000000005C6;
assign u[4'b1000] [07] = 64'h00000000000009C6;
assign v[4'b1000] [07] = 64'h0000000000000DC6;
assign X[4'b1000] [08] = 64'h0000000000000207;
assign Y[4'b1000] [08] = 64'h00000000000005C7;
assign u[4'b1000] [08] = 64'h00000000000009C7;
assign v[4'b1000] [08] = 64'h0000000000000DC7;
assign X[4'b1000] [09] = 64'h0000000000000208;
assign Y[4'b1000] [09] = 64'h00000000000005C8;
assign u[4'b1000] [09] = 64'h00000000000009C8;
assign v[4'b1000] [09] = 64'h0000000000000DC8;
assign X[4'b1000] [10] = 64'h0000000000000209;
assign Y[4'b1000] [10] = 64'h00000000000005C9;
assign u[4'b1000] [10] = 64'h00000000000009C9;
assign v[4'b1000] [10] = 64'h0000000000000DC9;
assign X[4'b1000] [11] = 64'h000000000000020A;
assign Y[4'b1000] [11] = 64'h00000000000005CA;
assign u[4'b1000] [11] = 64'h00000000000009CA;
assign v[4'b1000] [11] = 64'h0000000000000DCA;
assign X[4'b1000] [12] = 64'h000000000000020B;
assign Y[4'b1000] [12] = 64'h00000000000005CB;
assign u[4'b1000] [12] = 64'h00000000000009CB;
assign v[4'b1000] [12] = 64'h0000000000000DCB;
assign X[4'b1000] [13] = 64'h000000000000020C;
assign Y[4'b1000] [13] = 64'h00000000000005CC;
assign u[4'b1000] [13] = 64'h00000000000009CC;
assign v[4'b1000] [13] = 64'h0000000000000DCC;
assign X[4'b1000] [14] = 64'h000000000000020D;
assign Y[4'b1000] [14] = 64'h00000000000005CD;
assign u[4'b1000] [14] = 64'h00000000000009CD;
assign v[4'b1000] [14] = 64'h0000000000000DCD;
assign X[4'b1000] [15] = 64'h000000000000020E;
assign Y[4'b1000] [15] = 64'h00000000000005CE;
assign u[4'b1000] [15] = 64'h00000000000009CE;
assign v[4'b1000] [15] = 64'h0000000000000DCE;
assign X[4'b1000] [16] = 64'h000000000000020F;
assign Y[4'b1000] [16] = 64'h00000000000005CF;
assign u[4'b1000] [16] = 64'h00000000000009CF;
assign v[4'b1000] [16] = 64'h0000000000000DCF;
assign X[4'b1000] [17] = 64'h0000000000000210;
assign Y[4'b1000] [17] = 64'h00000000000005D0;
assign u[4'b1000] [17] = 64'h00000000000009D0;
assign v[4'b1000] [17] = 64'h0000000000000DD0;
assign X[4'b1000] [18] = 64'h0000000000000211;
assign Y[4'b1000] [18] = 64'h00000000000005D1;
assign u[4'b1000] [18] = 64'h00000000000009D1;
assign v[4'b1000] [18] = 64'h0000000000000DD1;
assign X[4'b1000] [19] = 64'h0000000000000212;
assign Y[4'b1000] [19] = 64'h00000000000005D2;
assign u[4'b1000] [19] = 64'h00000000000009D2;
assign v[4'b1000] [19] = 64'h0000000000000DD2;
assign X[4'b1000] [20] = 64'h0000000000000213;
assign Y[4'b1000] [20] = 64'h00000000000005D3;
assign u[4'b1000] [20] = 64'h00000000000009D3;
assign v[4'b1000] [20] = 64'h0000000000000DD3;
assign X[4'b1000] [21] = 64'h0000000000000214;
assign Y[4'b1000] [21] = 64'h00000000000005D4;
assign u[4'b1000] [21] = 64'h00000000000009D4;
assign v[4'b1000] [21] = 64'h0000000000000DD4;
assign X[4'b1000] [22] = 64'h0000000000000215;
assign Y[4'b1000] [22] = 64'h00000000000005D5;
assign u[4'b1000] [22] = 64'h00000000000009D5;
assign v[4'b1000] [22] = 64'h0000000000000DD5;
assign X[4'b1000] [23] = 64'h0000000000000216;
assign Y[4'b1000] [23] = 64'h00000000000005D6;
assign u[4'b1000] [23] = 64'h00000000000009D6;
assign v[4'b1000] [23] = 64'h0000000000000DD6;
assign X[4'b1000] [24] = 64'h0000000000000217;
assign Y[4'b1000] [24] = 64'h00000000000005D7;
assign u[4'b1000] [24] = 64'h00000000000009D7;
assign v[4'b1000] [24] = 64'h0000000000000DD7;
assign X[4'b1000] [25] = 64'h0000000000000218;
assign Y[4'b1000] [25] = 64'h00000000000005D8;
assign u[4'b1000] [25] = 64'h00000000000009D8;
assign v[4'b1000] [25] = 64'h0000000000000DD8;
assign X[4'b1000] [26] = 64'h0000000000000219;
assign Y[4'b1000] [26] = 64'h00000000000005D9;
assign u[4'b1000] [26] = 64'h00000000000009D9;
assign v[4'b1000] [26] = 64'h0000000000000DD9;
assign X[4'b1000] [27] = 64'h000000000000021A;
assign Y[4'b1000] [27] = 64'h00000000000005DA;
assign u[4'b1000] [27] = 64'h00000000000009DA;
assign v[4'b1000] [27] = 64'h0000000000000DDA;
assign X[4'b1000] [28] = 64'h000000000000021B;
assign Y[4'b1000] [28] = 64'h00000000000005DB;
assign u[4'b1000] [28] = 64'h00000000000009DB;
assign v[4'b1000] [28] = 64'h0000000000000DDB;
assign X[4'b1000] [29] = 64'h000000000000021C;
assign Y[4'b1000] [29] = 64'h00000000000005DC;
assign u[4'b1000] [29] = 64'h00000000000009DC;
assign v[4'b1000] [29] = 64'h0000000000000DDC;
assign X[4'b1000] [30] = 64'h000000000000021D;
assign Y[4'b1000] [30] = 64'h00000000000005DD;
assign u[4'b1000] [30] = 64'h00000000000009DD;
assign v[4'b1000] [30] = 64'h0000000000000DDD;
assign X[4'b1000] [31] = 64'h000000000000021E;
assign Y[4'b1000] [31] = 64'h00000000000005DE;
assign u[4'b1000] [31] = 64'h00000000000009DE;
assign v[4'b1000] [31] = 64'h0000000000000DDE;
assign X[4'b1000] [32] = 64'h000000000000021F;
assign Y[4'b1000] [32] = 64'h00000000000005DF;
assign u[4'b1000] [32] = 64'h00000000000009DF;
assign v[4'b1000] [32] = 64'h0000000000000DDF;
assign X[4'b1000] [33] = 64'h0000000000000220;
assign Y[4'b1000] [33] = 64'h00000000000005E0;
assign u[4'b1000] [33] = 64'h00000000000009E0;
assign v[4'b1000] [33] = 64'h0000000000000DE0;
assign X[4'b1000] [34] = 64'h0000000000000221;
assign Y[4'b1000] [34] = 64'h00000000000005E1;
assign u[4'b1000] [34] = 64'h00000000000009E1;
assign v[4'b1000] [34] = 64'h0000000000000DE1;
assign X[4'b1000] [35] = 64'h0000000000000222;
assign Y[4'b1000] [35] = 64'h00000000000005E2;
assign u[4'b1000] [35] = 64'h00000000000009E2;
assign v[4'b1000] [35] = 64'h0000000000000DE2;
assign X[4'b1000] [36] = 64'h0000000000000223;
assign Y[4'b1000] [36] = 64'h00000000000005E3;
assign u[4'b1000] [36] = 64'h00000000000009E3;
assign v[4'b1000] [36] = 64'h0000000000000DE3;
assign X[4'b1000] [37] = 64'h0000000000000224;
assign Y[4'b1000] [37] = 64'h00000000000005E4;
assign u[4'b1000] [37] = 64'h00000000000009E4;
assign v[4'b1000] [37] = 64'h0000000000000DE4;
assign X[4'b1000] [38] = 64'h0000000000000225;
assign Y[4'b1000] [38] = 64'h00000000000005E5;
assign u[4'b1000] [38] = 64'h00000000000009E5;
assign v[4'b1000] [38] = 64'h0000000000000DE5;
assign X[4'b1000] [39] = 64'h0000000000000226;
assign Y[4'b1000] [39] = 64'h00000000000005E6;
assign u[4'b1000] [39] = 64'h00000000000009E6;
assign v[4'b1000] [39] = 64'h0000000000000DE6;
assign X[4'b1000] [40] = 64'h0000000000000227;
assign Y[4'b1000] [40] = 64'h00000000000005E7;
assign u[4'b1000] [40] = 64'h00000000000009E7;
assign v[4'b1000] [40] = 64'h0000000000000DE7;
assign X[4'b1000] [41] = 64'h0000000000000228;
assign Y[4'b1000] [41] = 64'h00000000000005E8;
assign u[4'b1000] [41] = 64'h00000000000009E8;
assign v[4'b1000] [41] = 64'h0000000000000DE8;
assign X[4'b1000] [42] = 64'h0000000000000229;
assign Y[4'b1000] [42] = 64'h00000000000005E9;
assign u[4'b1000] [42] = 64'h00000000000009E9;
assign v[4'b1000] [42] = 64'h0000000000000DE9;
assign X[4'b1000] [43] = 64'h000000000000022A;
assign Y[4'b1000] [43] = 64'h00000000000005EA;
assign u[4'b1000] [43] = 64'h00000000000009EA;
assign v[4'b1000] [43] = 64'h0000000000000DEA;
assign X[4'b1000] [44] = 64'h000000000000022B;
assign Y[4'b1000] [44] = 64'h00000000000005EB;
assign u[4'b1000] [44] = 64'h00000000000009EB;
assign v[4'b1000] [44] = 64'h0000000000000DEB;
assign X[4'b1000] [45] = 64'h000000000000022C;
assign Y[4'b1000] [45] = 64'h00000000000005EC;
assign u[4'b1000] [45] = 64'h00000000000009EC;
assign v[4'b1000] [45] = 64'h0000000000000DEC;
assign X[4'b1000] [46] = 64'h000000000000022D;
assign Y[4'b1000] [46] = 64'h00000000000005ED;
assign u[4'b1000] [46] = 64'h00000000000009ED;
assign v[4'b1000] [46] = 64'h0000000000000DED;
assign X[4'b1000] [47] = 64'h000000000000022E;
assign Y[4'b1000] [47] = 64'h00000000000005EE;
assign u[4'b1000] [47] = 64'h00000000000009EE;
assign v[4'b1000] [47] = 64'h0000000000000DEE;
assign X[4'b1000] [48] = 64'h000000000000022F;
assign Y[4'b1000] [48] = 64'h00000000000005EF;
assign u[4'b1000] [48] = 64'h00000000000009EF;
assign v[4'b1000] [48] = 64'h0000000000000DEF;
assign X[4'b1000] [49] = 64'h0000000000000230;
assign Y[4'b1000] [49] = 64'h00000000000005F0;
assign u[4'b1000] [49] = 64'h00000000000009F0;
assign v[4'b1000] [49] = 64'h0000000000000DF0;
assign X[4'b1000] [50] = 64'h0000000000000231;
assign Y[4'b1000] [50] = 64'h00000000000005F1;
assign u[4'b1000] [50] = 64'h00000000000009F1;
assign v[4'b1000] [50] = 64'h0000000000000DF1;
assign X[4'b1000] [51] = 64'h0000000000000232;
assign Y[4'b1000] [51] = 64'h00000000000005F2;
assign u[4'b1000] [51] = 64'h00000000000009F2;
assign v[4'b1000] [51] = 64'h0000000000000DF2;
assign X[4'b1000] [52] = 64'h0000000000000233;
assign Y[4'b1000] [52] = 64'h00000000000005F3;
assign u[4'b1000] [52] = 64'h00000000000009F3;
assign v[4'b1000] [52] = 64'h0000000000000DF3;
assign X[4'b1000] [53] = 64'h0000000000000234;
assign Y[4'b1000] [53] = 64'h00000000000005F4;
assign u[4'b1000] [53] = 64'h00000000000009F4;
assign v[4'b1000] [53] = 64'h0000000000000DF4;
assign X[4'b1000] [54] = 64'h0000000000000235;
assign Y[4'b1000] [54] = 64'h00000000000005F5;
assign u[4'b1000] [54] = 64'h00000000000009F5;
assign v[4'b1000] [54] = 64'h0000000000000DF5;
assign X[4'b1000] [55] = 64'h0000000000000236;
assign Y[4'b1000] [55] = 64'h00000000000005F6;
assign u[4'b1000] [55] = 64'h00000000000009F6;
assign v[4'b1000] [55] = 64'h0000000000000DF6;
assign X[4'b1000] [56] = 64'h0000000000000237;
assign Y[4'b1000] [56] = 64'h00000000000005F7;
assign u[4'b1000] [56] = 64'h00000000000009F7;
assign v[4'b1000] [56] = 64'h0000000000000DF7;
assign X[4'b1000] [57] = 64'h0000000000000238;
assign Y[4'b1000] [57] = 64'h00000000000005F8;
assign u[4'b1000] [57] = 64'h00000000000009F8;
assign v[4'b1000] [57] = 64'h0000000000000DF8;
assign X[4'b1000] [58] = 64'h0000000000000239;
assign Y[4'b1000] [58] = 64'h00000000000005F9;
assign u[4'b1000] [58] = 64'h00000000000009F9;
assign v[4'b1000] [58] = 64'h0000000000000DF9;
assign X[4'b1000] [59] = 64'h000000000000023A;
assign Y[4'b1000] [59] = 64'h00000000000005FA;
assign u[4'b1000] [59] = 64'h00000000000009FA;
assign v[4'b1000] [59] = 64'h0000000000000DFA;
assign X[4'b1000] [60] = 64'h000000000000023B;
assign Y[4'b1000] [60] = 64'h00000000000005FB;
assign u[4'b1000] [60] = 64'h00000000000009FB;
assign v[4'b1000] [60] = 64'h0000000000000DFB;
assign X[4'b1000] [61] = 64'h000000000000023C;
assign Y[4'b1000] [61] = 64'h00000000000005FC;
assign u[4'b1000] [61] = 64'h00000000000009FC;
assign v[4'b1000] [61] = 64'h0000000000000DFC;
assign X[4'b1000] [62] = 64'h000000000000023D;
assign Y[4'b1000] [62] = 64'h00000000000005FD;
assign u[4'b1000] [62] = 64'h00000000000009FD;
assign v[4'b1000] [62] = 64'h0000000000000DFD;
assign X[4'b1000] [63] = 64'h000000000000023E;
assign Y[4'b1000] [63] = 64'h00000000000005FE;
assign u[4'b1000] [63] = 64'h00000000000009FE;
assign v[4'b1000] [63] = 64'h0000000000000DFE;
assign X[4'b1000] [64] = 64'h000000000000023F;
assign Y[4'b1000] [64] = 64'h00000000000005FF;
assign u[4'b1000] [64] = 64'h00000000000009FF;
assign v[4'b1000] [64] = 64'h0000000000000DFF;
assign X[4'b1001] [01] = 64'h0000000000000240;
assign Y[4'b1001] [01] = 64'h0000000000000600;
assign u[4'b1001] [01] = 64'h0000000000000A00;
assign v[4'b1001] [01] = 64'h0000000000000E00;
assign X[4'b1001] [02] = 64'h0000000000000241;
assign Y[4'b1001] [02] = 64'h0000000000000601;
assign u[4'b1001] [02] = 64'h0000000000000A01;
assign v[4'b1001] [02] = 64'h0000000000000E01;
assign X[4'b1001] [03] = 64'h0000000000000242;
assign Y[4'b1001] [03] = 64'h0000000000000602;
assign u[4'b1001] [03] = 64'h0000000000000A02;
assign v[4'b1001] [03] = 64'h0000000000000E02;
assign X[4'b1001] [04] = 64'h0000000000000243;
assign Y[4'b1001] [04] = 64'h0000000000000603;
assign u[4'b1001] [04] = 64'h0000000000000A03;
assign v[4'b1001] [04] = 64'h0000000000000E03;
assign X[4'b1001] [05] = 64'h0000000000000244;
assign Y[4'b1001] [05] = 64'h0000000000000604;
assign u[4'b1001] [05] = 64'h0000000000000A04;
assign v[4'b1001] [05] = 64'h0000000000000E04;
assign X[4'b1001] [06] = 64'h0000000000000245;
assign Y[4'b1001] [06] = 64'h0000000000000605;
assign u[4'b1001] [06] = 64'h0000000000000A05;
assign v[4'b1001] [06] = 64'h0000000000000E05;
assign X[4'b1001] [07] = 64'h0000000000000246;
assign Y[4'b1001] [07] = 64'h0000000000000606;
assign u[4'b1001] [07] = 64'h0000000000000A06;
assign v[4'b1001] [07] = 64'h0000000000000E06;
assign X[4'b1001] [08] = 64'h0000000000000247;
assign Y[4'b1001] [08] = 64'h0000000000000607;
assign u[4'b1001] [08] = 64'h0000000000000A07;
assign v[4'b1001] [08] = 64'h0000000000000E07;
assign X[4'b1001] [09] = 64'h0000000000000248;
assign Y[4'b1001] [09] = 64'h0000000000000608;
assign u[4'b1001] [09] = 64'h0000000000000A08;
assign v[4'b1001] [09] = 64'h0000000000000E08;
assign X[4'b1001] [10] = 64'h0000000000000249;
assign Y[4'b1001] [10] = 64'h0000000000000609;
assign u[4'b1001] [10] = 64'h0000000000000A09;
assign v[4'b1001] [10] = 64'h0000000000000E09;
assign X[4'b1001] [11] = 64'h000000000000024A;
assign Y[4'b1001] [11] = 64'h000000000000060A;
assign u[4'b1001] [11] = 64'h0000000000000A0A;
assign v[4'b1001] [11] = 64'h0000000000000E0A;
assign X[4'b1001] [12] = 64'h000000000000024B;
assign Y[4'b1001] [12] = 64'h000000000000060B;
assign u[4'b1001] [12] = 64'h0000000000000A0B;
assign v[4'b1001] [12] = 64'h0000000000000E0B;
assign X[4'b1001] [13] = 64'h000000000000024C;
assign Y[4'b1001] [13] = 64'h000000000000060C;
assign u[4'b1001] [13] = 64'h0000000000000A0C;
assign v[4'b1001] [13] = 64'h0000000000000E0C;
assign X[4'b1001] [14] = 64'h000000000000024D;
assign Y[4'b1001] [14] = 64'h000000000000060D;
assign u[4'b1001] [14] = 64'h0000000000000A0D;
assign v[4'b1001] [14] = 64'h0000000000000E0D;
assign X[4'b1001] [15] = 64'h000000000000024E;
assign Y[4'b1001] [15] = 64'h000000000000060E;
assign u[4'b1001] [15] = 64'h0000000000000A0E;
assign v[4'b1001] [15] = 64'h0000000000000E0E;
assign X[4'b1001] [16] = 64'h000000000000024F;
assign Y[4'b1001] [16] = 64'h000000000000060F;
assign u[4'b1001] [16] = 64'h0000000000000A0F;
assign v[4'b1001] [16] = 64'h0000000000000E0F;
assign X[4'b1001] [17] = 64'h0000000000000250;
assign Y[4'b1001] [17] = 64'h0000000000000610;
assign u[4'b1001] [17] = 64'h0000000000000A10;
assign v[4'b1001] [17] = 64'h0000000000000E10;
assign X[4'b1001] [18] = 64'h0000000000000251;
assign Y[4'b1001] [18] = 64'h0000000000000611;
assign u[4'b1001] [18] = 64'h0000000000000A11;
assign v[4'b1001] [18] = 64'h0000000000000E11;
assign X[4'b1001] [19] = 64'h0000000000000252;
assign Y[4'b1001] [19] = 64'h0000000000000612;
assign u[4'b1001] [19] = 64'h0000000000000A12;
assign v[4'b1001] [19] = 64'h0000000000000E12;
assign X[4'b1001] [20] = 64'h0000000000000253;
assign Y[4'b1001] [20] = 64'h0000000000000613;
assign u[4'b1001] [20] = 64'h0000000000000A13;
assign v[4'b1001] [20] = 64'h0000000000000E13;
assign X[4'b1001] [21] = 64'h0000000000000254;
assign Y[4'b1001] [21] = 64'h0000000000000614;
assign u[4'b1001] [21] = 64'h0000000000000A14;
assign v[4'b1001] [21] = 64'h0000000000000E14;
assign X[4'b1001] [22] = 64'h0000000000000255;
assign Y[4'b1001] [22] = 64'h0000000000000615;
assign u[4'b1001] [22] = 64'h0000000000000A15;
assign v[4'b1001] [22] = 64'h0000000000000E15;
assign X[4'b1001] [23] = 64'h0000000000000256;
assign Y[4'b1001] [23] = 64'h0000000000000616;
assign u[4'b1001] [23] = 64'h0000000000000A16;
assign v[4'b1001] [23] = 64'h0000000000000E16;
assign X[4'b1001] [24] = 64'h0000000000000257;
assign Y[4'b1001] [24] = 64'h0000000000000617;
assign u[4'b1001] [24] = 64'h0000000000000A17;
assign v[4'b1001] [24] = 64'h0000000000000E17;
assign X[4'b1001] [25] = 64'h0000000000000258;
assign Y[4'b1001] [25] = 64'h0000000000000618;
assign u[4'b1001] [25] = 64'h0000000000000A18;
assign v[4'b1001] [25] = 64'h0000000000000E18;
assign X[4'b1001] [26] = 64'h0000000000000259;
assign Y[4'b1001] [26] = 64'h0000000000000619;
assign u[4'b1001] [26] = 64'h0000000000000A19;
assign v[4'b1001] [26] = 64'h0000000000000E19;
assign X[4'b1001] [27] = 64'h000000000000025A;
assign Y[4'b1001] [27] = 64'h000000000000061A;
assign u[4'b1001] [27] = 64'h0000000000000A1A;
assign v[4'b1001] [27] = 64'h0000000000000E1A;
assign X[4'b1001] [28] = 64'h000000000000025B;
assign Y[4'b1001] [28] = 64'h000000000000061B;
assign u[4'b1001] [28] = 64'h0000000000000A1B;
assign v[4'b1001] [28] = 64'h0000000000000E1B;
assign X[4'b1001] [29] = 64'h000000000000025C;
assign Y[4'b1001] [29] = 64'h000000000000061C;
assign u[4'b1001] [29] = 64'h0000000000000A1C;
assign v[4'b1001] [29] = 64'h0000000000000E1C;
assign X[4'b1001] [30] = 64'h000000000000025D;
assign Y[4'b1001] [30] = 64'h000000000000061D;
assign u[4'b1001] [30] = 64'h0000000000000A1D;
assign v[4'b1001] [30] = 64'h0000000000000E1D;
assign X[4'b1001] [31] = 64'h000000000000025E;
assign Y[4'b1001] [31] = 64'h000000000000061E;
assign u[4'b1001] [31] = 64'h0000000000000A1E;
assign v[4'b1001] [31] = 64'h0000000000000E1E;
assign X[4'b1001] [32] = 64'h000000000000025F;
assign Y[4'b1001] [32] = 64'h000000000000061F;
assign u[4'b1001] [32] = 64'h0000000000000A1F;
assign v[4'b1001] [32] = 64'h0000000000000E1F;
assign X[4'b1001] [33] = 64'h0000000000000260;
assign Y[4'b1001] [33] = 64'h0000000000000620;
assign u[4'b1001] [33] = 64'h0000000000000A20;
assign v[4'b1001] [33] = 64'h0000000000000E20;
assign X[4'b1001] [34] = 64'h0000000000000261;
assign Y[4'b1001] [34] = 64'h0000000000000621;
assign u[4'b1001] [34] = 64'h0000000000000A21;
assign v[4'b1001] [34] = 64'h0000000000000E21;
assign X[4'b1001] [35] = 64'h0000000000000262;
assign Y[4'b1001] [35] = 64'h0000000000000622;
assign u[4'b1001] [35] = 64'h0000000000000A22;
assign v[4'b1001] [35] = 64'h0000000000000E22;
assign X[4'b1001] [36] = 64'h0000000000000263;
assign Y[4'b1001] [36] = 64'h0000000000000623;
assign u[4'b1001] [36] = 64'h0000000000000A23;
assign v[4'b1001] [36] = 64'h0000000000000E23;
assign X[4'b1001] [37] = 64'h0000000000000264;
assign Y[4'b1001] [37] = 64'h0000000000000624;
assign u[4'b1001] [37] = 64'h0000000000000A24;
assign v[4'b1001] [37] = 64'h0000000000000E24;
assign X[4'b1001] [38] = 64'h0000000000000265;
assign Y[4'b1001] [38] = 64'h0000000000000625;
assign u[4'b1001] [38] = 64'h0000000000000A25;
assign v[4'b1001] [38] = 64'h0000000000000E25;
assign X[4'b1001] [39] = 64'h0000000000000266;
assign Y[4'b1001] [39] = 64'h0000000000000626;
assign u[4'b1001] [39] = 64'h0000000000000A26;
assign v[4'b1001] [39] = 64'h0000000000000E26;
assign X[4'b1001] [40] = 64'h0000000000000267;
assign Y[4'b1001] [40] = 64'h0000000000000627;
assign u[4'b1001] [40] = 64'h0000000000000A27;
assign v[4'b1001] [40] = 64'h0000000000000E27;
assign X[4'b1001] [41] = 64'h0000000000000268;
assign Y[4'b1001] [41] = 64'h0000000000000628;
assign u[4'b1001] [41] = 64'h0000000000000A28;
assign v[4'b1001] [41] = 64'h0000000000000E28;
assign X[4'b1001] [42] = 64'h0000000000000269;
assign Y[4'b1001] [42] = 64'h0000000000000629;
assign u[4'b1001] [42] = 64'h0000000000000A29;
assign v[4'b1001] [42] = 64'h0000000000000E29;
assign X[4'b1001] [43] = 64'h000000000000026A;
assign Y[4'b1001] [43] = 64'h000000000000062A;
assign u[4'b1001] [43] = 64'h0000000000000A2A;
assign v[4'b1001] [43] = 64'h0000000000000E2A;
assign X[4'b1001] [44] = 64'h000000000000026B;
assign Y[4'b1001] [44] = 64'h000000000000062B;
assign u[4'b1001] [44] = 64'h0000000000000A2B;
assign v[4'b1001] [44] = 64'h0000000000000E2B;
assign X[4'b1001] [45] = 64'h000000000000026C;
assign Y[4'b1001] [45] = 64'h000000000000062C;
assign u[4'b1001] [45] = 64'h0000000000000A2C;
assign v[4'b1001] [45] = 64'h0000000000000E2C;
assign X[4'b1001] [46] = 64'h000000000000026D;
assign Y[4'b1001] [46] = 64'h000000000000062D;
assign u[4'b1001] [46] = 64'h0000000000000A2D;
assign v[4'b1001] [46] = 64'h0000000000000E2D;
assign X[4'b1001] [47] = 64'h000000000000026E;
assign Y[4'b1001] [47] = 64'h000000000000062E;
assign u[4'b1001] [47] = 64'h0000000000000A2E;
assign v[4'b1001] [47] = 64'h0000000000000E2E;
assign X[4'b1001] [48] = 64'h000000000000026F;
assign Y[4'b1001] [48] = 64'h000000000000062F;
assign u[4'b1001] [48] = 64'h0000000000000A2F;
assign v[4'b1001] [48] = 64'h0000000000000E2F;
assign X[4'b1001] [49] = 64'h0000000000000270;
assign Y[4'b1001] [49] = 64'h0000000000000630;
assign u[4'b1001] [49] = 64'h0000000000000A30;
assign v[4'b1001] [49] = 64'h0000000000000E30;
assign X[4'b1001] [50] = 64'h0000000000000271;
assign Y[4'b1001] [50] = 64'h0000000000000631;
assign u[4'b1001] [50] = 64'h0000000000000A31;
assign v[4'b1001] [50] = 64'h0000000000000E31;
assign X[4'b1001] [51] = 64'h0000000000000272;
assign Y[4'b1001] [51] = 64'h0000000000000632;
assign u[4'b1001] [51] = 64'h0000000000000A32;
assign v[4'b1001] [51] = 64'h0000000000000E32;
assign X[4'b1001] [52] = 64'h0000000000000273;
assign Y[4'b1001] [52] = 64'h0000000000000633;
assign u[4'b1001] [52] = 64'h0000000000000A33;
assign v[4'b1001] [52] = 64'h0000000000000E33;
assign X[4'b1001] [53] = 64'h0000000000000274;
assign Y[4'b1001] [53] = 64'h0000000000000634;
assign u[4'b1001] [53] = 64'h0000000000000A34;
assign v[4'b1001] [53] = 64'h0000000000000E34;
assign X[4'b1001] [54] = 64'h0000000000000275;
assign Y[4'b1001] [54] = 64'h0000000000000635;
assign u[4'b1001] [54] = 64'h0000000000000A35;
assign v[4'b1001] [54] = 64'h0000000000000E35;
assign X[4'b1001] [55] = 64'h0000000000000276;
assign Y[4'b1001] [55] = 64'h0000000000000636;
assign u[4'b1001] [55] = 64'h0000000000000A36;
assign v[4'b1001] [55] = 64'h0000000000000E36;
assign X[4'b1001] [56] = 64'h0000000000000277;
assign Y[4'b1001] [56] = 64'h0000000000000637;
assign u[4'b1001] [56] = 64'h0000000000000A37;
assign v[4'b1001] [56] = 64'h0000000000000E37;
assign X[4'b1001] [57] = 64'h0000000000000278;
assign Y[4'b1001] [57] = 64'h0000000000000638;
assign u[4'b1001] [57] = 64'h0000000000000A38;
assign v[4'b1001] [57] = 64'h0000000000000E38;
assign X[4'b1001] [58] = 64'h0000000000000279;
assign Y[4'b1001] [58] = 64'h0000000000000639;
assign u[4'b1001] [58] = 64'h0000000000000A39;
assign v[4'b1001] [58] = 64'h0000000000000E39;
assign X[4'b1001] [59] = 64'h000000000000027A;
assign Y[4'b1001] [59] = 64'h000000000000063A;
assign u[4'b1001] [59] = 64'h0000000000000A3A;
assign v[4'b1001] [59] = 64'h0000000000000E3A;
assign X[4'b1001] [60] = 64'h000000000000027B;
assign Y[4'b1001] [60] = 64'h000000000000063B;
assign u[4'b1001] [60] = 64'h0000000000000A3B;
assign v[4'b1001] [60] = 64'h0000000000000E3B;
assign X[4'b1001] [61] = 64'h000000000000027C;
assign Y[4'b1001] [61] = 64'h000000000000063C;
assign u[4'b1001] [61] = 64'h0000000000000A3C;
assign v[4'b1001] [61] = 64'h0000000000000E3C;
assign X[4'b1001] [62] = 64'h000000000000027D;
assign Y[4'b1001] [62] = 64'h000000000000063D;
assign u[4'b1001] [62] = 64'h0000000000000A3D;
assign v[4'b1001] [62] = 64'h0000000000000E3D;
assign X[4'b1001] [63] = 64'h000000000000027E;
assign Y[4'b1001] [63] = 64'h000000000000063E;
assign u[4'b1001] [63] = 64'h0000000000000A3E;
assign v[4'b1001] [63] = 64'h0000000000000E3E;
assign X[4'b1001] [64] = 64'h000000000000027F;
assign Y[4'b1001] [64] = 64'h000000000000063F;
assign u[4'b1001] [64] = 64'h0000000000000A3F;
assign v[4'b1001] [64] = 64'h0000000000000E3F;
assign X[4'b1010] [01] = 64'h0000000000000280;
assign Y[4'b1010] [01] = 64'h0000000000000640;
assign u[4'b1010] [01] = 64'h0000000000000A40;
assign v[4'b1010] [01] = 64'h0000000000000E40;
assign X[4'b1010] [02] = 64'h0000000000000281;
assign Y[4'b1010] [02] = 64'h0000000000000641;
assign u[4'b1010] [02] = 64'h0000000000000A41;
assign v[4'b1010] [02] = 64'h0000000000000E41;
assign X[4'b1010] [03] = 64'h0000000000000282;
assign Y[4'b1010] [03] = 64'h0000000000000642;
assign u[4'b1010] [03] = 64'h0000000000000A42;
assign v[4'b1010] [03] = 64'h0000000000000E42;
assign X[4'b1010] [04] = 64'h0000000000000283;
assign Y[4'b1010] [04] = 64'h0000000000000643;
assign u[4'b1010] [04] = 64'h0000000000000A43;
assign v[4'b1010] [04] = 64'h0000000000000E43;
assign X[4'b1010] [05] = 64'h0000000000000284;
assign Y[4'b1010] [05] = 64'h0000000000000644;
assign u[4'b1010] [05] = 64'h0000000000000A44;
assign v[4'b1010] [05] = 64'h0000000000000E44;
assign X[4'b1010] [06] = 64'h0000000000000285;
assign Y[4'b1010] [06] = 64'h0000000000000645;
assign u[4'b1010] [06] = 64'h0000000000000A45;
assign v[4'b1010] [06] = 64'h0000000000000E45;
assign X[4'b1010] [07] = 64'h0000000000000286;
assign Y[4'b1010] [07] = 64'h0000000000000646;
assign u[4'b1010] [07] = 64'h0000000000000A46;
assign v[4'b1010] [07] = 64'h0000000000000E46;
assign X[4'b1010] [08] = 64'h0000000000000287;
assign Y[4'b1010] [08] = 64'h0000000000000647;
assign u[4'b1010] [08] = 64'h0000000000000A47;
assign v[4'b1010] [08] = 64'h0000000000000E47;
assign X[4'b1010] [09] = 64'h0000000000000288;
assign Y[4'b1010] [09] = 64'h0000000000000648;
assign u[4'b1010] [09] = 64'h0000000000000A48;
assign v[4'b1010] [09] = 64'h0000000000000E48;
assign X[4'b1010] [10] = 64'h0000000000000289;
assign Y[4'b1010] [10] = 64'h0000000000000649;
assign u[4'b1010] [10] = 64'h0000000000000A49;
assign v[4'b1010] [10] = 64'h0000000000000E49;
assign X[4'b1010] [11] = 64'h000000000000028A;
assign Y[4'b1010] [11] = 64'h000000000000064A;
assign u[4'b1010] [11] = 64'h0000000000000A4A;
assign v[4'b1010] [11] = 64'h0000000000000E4A;
assign X[4'b1010] [12] = 64'h000000000000028B;
assign Y[4'b1010] [12] = 64'h000000000000064B;
assign u[4'b1010] [12] = 64'h0000000000000A4B;
assign v[4'b1010] [12] = 64'h0000000000000E4B;
assign X[4'b1010] [13] = 64'h000000000000028C;
assign Y[4'b1010] [13] = 64'h000000000000064C;
assign u[4'b1010] [13] = 64'h0000000000000A4C;
assign v[4'b1010] [13] = 64'h0000000000000E4C;
assign X[4'b1010] [14] = 64'h000000000000028D;
assign Y[4'b1010] [14] = 64'h000000000000064D;
assign u[4'b1010] [14] = 64'h0000000000000A4D;
assign v[4'b1010] [14] = 64'h0000000000000E4D;
assign X[4'b1010] [15] = 64'h000000000000028E;
assign Y[4'b1010] [15] = 64'h000000000000064E;
assign u[4'b1010] [15] = 64'h0000000000000A4E;
assign v[4'b1010] [15] = 64'h0000000000000E4E;
assign X[4'b1010] [16] = 64'h000000000000028F;
assign Y[4'b1010] [16] = 64'h000000000000064F;
assign u[4'b1010] [16] = 64'h0000000000000A4F;
assign v[4'b1010] [16] = 64'h0000000000000E4F;
assign X[4'b1010] [17] = 64'h0000000000000290;
assign Y[4'b1010] [17] = 64'h0000000000000650;
assign u[4'b1010] [17] = 64'h0000000000000A50;
assign v[4'b1010] [17] = 64'h0000000000000E50;
assign X[4'b1010] [18] = 64'h0000000000000291;
assign Y[4'b1010] [18] = 64'h0000000000000651;
assign u[4'b1010] [18] = 64'h0000000000000A51;
assign v[4'b1010] [18] = 64'h0000000000000E51;
assign X[4'b1010] [19] = 64'h0000000000000292;
assign Y[4'b1010] [19] = 64'h0000000000000652;
assign u[4'b1010] [19] = 64'h0000000000000A52;
assign v[4'b1010] [19] = 64'h0000000000000E52;
assign X[4'b1010] [20] = 64'h0000000000000293;
assign Y[4'b1010] [20] = 64'h0000000000000653;
assign u[4'b1010] [20] = 64'h0000000000000A53;
assign v[4'b1010] [20] = 64'h0000000000000E53;
assign X[4'b1010] [21] = 64'h0000000000000294;
assign Y[4'b1010] [21] = 64'h0000000000000654;
assign u[4'b1010] [21] = 64'h0000000000000A54;
assign v[4'b1010] [21] = 64'h0000000000000E54;
assign X[4'b1010] [22] = 64'h0000000000000295;
assign Y[4'b1010] [22] = 64'h0000000000000655;
assign u[4'b1010] [22] = 64'h0000000000000A55;
assign v[4'b1010] [22] = 64'h0000000000000E55;
assign X[4'b1010] [23] = 64'h0000000000000296;
assign Y[4'b1010] [23] = 64'h0000000000000656;
assign u[4'b1010] [23] = 64'h0000000000000A56;
assign v[4'b1010] [23] = 64'h0000000000000E56;
assign X[4'b1010] [24] = 64'h0000000000000297;
assign Y[4'b1010] [24] = 64'h0000000000000657;
assign u[4'b1010] [24] = 64'h0000000000000A57;
assign v[4'b1010] [24] = 64'h0000000000000E57;
assign X[4'b1010] [25] = 64'h0000000000000298;
assign Y[4'b1010] [25] = 64'h0000000000000658;
assign u[4'b1010] [25] = 64'h0000000000000A58;
assign v[4'b1010] [25] = 64'h0000000000000E58;
assign X[4'b1010] [26] = 64'h0000000000000299;
assign Y[4'b1010] [26] = 64'h0000000000000659;
assign u[4'b1010] [26] = 64'h0000000000000A59;
assign v[4'b1010] [26] = 64'h0000000000000E59;
assign X[4'b1010] [27] = 64'h000000000000029A;
assign Y[4'b1010] [27] = 64'h000000000000065A;
assign u[4'b1010] [27] = 64'h0000000000000A5A;
assign v[4'b1010] [27] = 64'h0000000000000E5A;
assign X[4'b1010] [28] = 64'h000000000000029B;
assign Y[4'b1010] [28] = 64'h000000000000065B;
assign u[4'b1010] [28] = 64'h0000000000000A5B;
assign v[4'b1010] [28] = 64'h0000000000000E5B;
assign X[4'b1010] [29] = 64'h000000000000029C;
assign Y[4'b1010] [29] = 64'h000000000000065C;
assign u[4'b1010] [29] = 64'h0000000000000A5C;
assign v[4'b1010] [29] = 64'h0000000000000E5C;
assign X[4'b1010] [30] = 64'h000000000000029D;
assign Y[4'b1010] [30] = 64'h000000000000065D;
assign u[4'b1010] [30] = 64'h0000000000000A5D;
assign v[4'b1010] [30] = 64'h0000000000000E5D;
assign X[4'b1010] [31] = 64'h000000000000029E;
assign Y[4'b1010] [31] = 64'h000000000000065E;
assign u[4'b1010] [31] = 64'h0000000000000A5E;
assign v[4'b1010] [31] = 64'h0000000000000E5E;
assign X[4'b1010] [32] = 64'h000000000000029F;
assign Y[4'b1010] [32] = 64'h000000000000065F;
assign u[4'b1010] [32] = 64'h0000000000000A5F;
assign v[4'b1010] [32] = 64'h0000000000000E5F;
assign X[4'b1010] [33] = 64'h00000000000002A0;
assign Y[4'b1010] [33] = 64'h0000000000000660;
assign u[4'b1010] [33] = 64'h0000000000000A60;
assign v[4'b1010] [33] = 64'h0000000000000E60;
assign X[4'b1010] [34] = 64'h00000000000002A1;
assign Y[4'b1010] [34] = 64'h0000000000000661;
assign u[4'b1010] [34] = 64'h0000000000000A61;
assign v[4'b1010] [34] = 64'h0000000000000E61;
assign X[4'b1010] [35] = 64'h00000000000002A2;
assign Y[4'b1010] [35] = 64'h0000000000000662;
assign u[4'b1010] [35] = 64'h0000000000000A62;
assign v[4'b1010] [35] = 64'h0000000000000E62;
assign X[4'b1010] [36] = 64'h00000000000002A3;
assign Y[4'b1010] [36] = 64'h0000000000000663;
assign u[4'b1010] [36] = 64'h0000000000000A63;
assign v[4'b1010] [36] = 64'h0000000000000E63;
assign X[4'b1010] [37] = 64'h00000000000002A4;
assign Y[4'b1010] [37] = 64'h0000000000000664;
assign u[4'b1010] [37] = 64'h0000000000000A64;
assign v[4'b1010] [37] = 64'h0000000000000E64;
assign X[4'b1010] [38] = 64'h00000000000002A5;
assign Y[4'b1010] [38] = 64'h0000000000000665;
assign u[4'b1010] [38] = 64'h0000000000000A65;
assign v[4'b1010] [38] = 64'h0000000000000E65;
assign X[4'b1010] [39] = 64'h00000000000002A6;
assign Y[4'b1010] [39] = 64'h0000000000000666;
assign u[4'b1010] [39] = 64'h0000000000000A66;
assign v[4'b1010] [39] = 64'h0000000000000E66;
assign X[4'b1010] [40] = 64'h00000000000002A7;
assign Y[4'b1010] [40] = 64'h0000000000000667;
assign u[4'b1010] [40] = 64'h0000000000000A67;
assign v[4'b1010] [40] = 64'h0000000000000E67;
assign X[4'b1010] [41] = 64'h00000000000002A8;
assign Y[4'b1010] [41] = 64'h0000000000000668;
assign u[4'b1010] [41] = 64'h0000000000000A68;
assign v[4'b1010] [41] = 64'h0000000000000E68;
assign X[4'b1010] [42] = 64'h00000000000002A9;
assign Y[4'b1010] [42] = 64'h0000000000000669;
assign u[4'b1010] [42] = 64'h0000000000000A69;
assign v[4'b1010] [42] = 64'h0000000000000E69;
assign X[4'b1010] [43] = 64'h00000000000002AA;
assign Y[4'b1010] [43] = 64'h000000000000066A;
assign u[4'b1010] [43] = 64'h0000000000000A6A;
assign v[4'b1010] [43] = 64'h0000000000000E6A;
assign X[4'b1010] [44] = 64'h00000000000002AB;
assign Y[4'b1010] [44] = 64'h000000000000066B;
assign u[4'b1010] [44] = 64'h0000000000000A6B;
assign v[4'b1010] [44] = 64'h0000000000000E6B;
assign X[4'b1010] [45] = 64'h00000000000002AC;
assign Y[4'b1010] [45] = 64'h000000000000066C;
assign u[4'b1010] [45] = 64'h0000000000000A6C;
assign v[4'b1010] [45] = 64'h0000000000000E6C;
assign X[4'b1010] [46] = 64'h00000000000002AD;
assign Y[4'b1010] [46] = 64'h000000000000066D;
assign u[4'b1010] [46] = 64'h0000000000000A6D;
assign v[4'b1010] [46] = 64'h0000000000000E6D;
assign X[4'b1010] [47] = 64'h00000000000002AE;
assign Y[4'b1010] [47] = 64'h000000000000066E;
assign u[4'b1010] [47] = 64'h0000000000000A6E;
assign v[4'b1010] [47] = 64'h0000000000000E6E;
assign X[4'b1010] [48] = 64'h00000000000002AF;
assign Y[4'b1010] [48] = 64'h000000000000066F;
assign u[4'b1010] [48] = 64'h0000000000000A6F;
assign v[4'b1010] [48] = 64'h0000000000000E6F;
assign X[4'b1010] [49] = 64'h00000000000002B0;
assign Y[4'b1010] [49] = 64'h0000000000000670;
assign u[4'b1010] [49] = 64'h0000000000000A70;
assign v[4'b1010] [49] = 64'h0000000000000E70;
assign X[4'b1010] [50] = 64'h00000000000002B1;
assign Y[4'b1010] [50] = 64'h0000000000000671;
assign u[4'b1010] [50] = 64'h0000000000000A71;
assign v[4'b1010] [50] = 64'h0000000000000E71;
assign X[4'b1010] [51] = 64'h00000000000002B2;
assign Y[4'b1010] [51] = 64'h0000000000000672;
assign u[4'b1010] [51] = 64'h0000000000000A72;
assign v[4'b1010] [51] = 64'h0000000000000E72;
assign X[4'b1010] [52] = 64'h00000000000002B3;
assign Y[4'b1010] [52] = 64'h0000000000000673;
assign u[4'b1010] [52] = 64'h0000000000000A73;
assign v[4'b1010] [52] = 64'h0000000000000E73;
assign X[4'b1010] [53] = 64'h00000000000002B4;
assign Y[4'b1010] [53] = 64'h0000000000000674;
assign u[4'b1010] [53] = 64'h0000000000000A74;
assign v[4'b1010] [53] = 64'h0000000000000E74;
assign X[4'b1010] [54] = 64'h00000000000002B5;
assign Y[4'b1010] [54] = 64'h0000000000000675;
assign u[4'b1010] [54] = 64'h0000000000000A75;
assign v[4'b1010] [54] = 64'h0000000000000E75;
assign X[4'b1010] [55] = 64'h00000000000002B6;
assign Y[4'b1010] [55] = 64'h0000000000000676;
assign u[4'b1010] [55] = 64'h0000000000000A76;
assign v[4'b1010] [55] = 64'h0000000000000E76;
assign X[4'b1010] [56] = 64'h00000000000002B7;
assign Y[4'b1010] [56] = 64'h0000000000000677;
assign u[4'b1010] [56] = 64'h0000000000000A77;
assign v[4'b1010] [56] = 64'h0000000000000E77;
assign X[4'b1010] [57] = 64'h00000000000002B8;
assign Y[4'b1010] [57] = 64'h0000000000000678;
assign u[4'b1010] [57] = 64'h0000000000000A78;
assign v[4'b1010] [57] = 64'h0000000000000E78;
assign X[4'b1010] [58] = 64'h00000000000002B9;
assign Y[4'b1010] [58] = 64'h0000000000000679;
assign u[4'b1010] [58] = 64'h0000000000000A79;
assign v[4'b1010] [58] = 64'h0000000000000E79;
assign X[4'b1010] [59] = 64'h00000000000002BA;
assign Y[4'b1010] [59] = 64'h000000000000067A;
assign u[4'b1010] [59] = 64'h0000000000000A7A;
assign v[4'b1010] [59] = 64'h0000000000000E7A;
assign X[4'b1010] [60] = 64'h00000000000002BB;
assign Y[4'b1010] [60] = 64'h000000000000067B;
assign u[4'b1010] [60] = 64'h0000000000000A7B;
assign v[4'b1010] [60] = 64'h0000000000000E7B;
assign X[4'b1010] [61] = 64'h00000000000002BC;
assign Y[4'b1010] [61] = 64'h000000000000067C;
assign u[4'b1010] [61] = 64'h0000000000000A7C;
assign v[4'b1010] [61] = 64'h0000000000000E7C;
assign X[4'b1010] [62] = 64'h00000000000002BD;
assign Y[4'b1010] [62] = 64'h000000000000067D;
assign u[4'b1010] [62] = 64'h0000000000000A7D;
assign v[4'b1010] [62] = 64'h0000000000000E7D;
assign X[4'b1010] [63] = 64'h00000000000002BE;
assign Y[4'b1010] [63] = 64'h000000000000067E;
assign u[4'b1010] [63] = 64'h0000000000000A7E;
assign v[4'b1010] [63] = 64'h0000000000000E7E;
assign X[4'b1010] [64] = 64'h00000000000002BF;
assign Y[4'b1010] [64] = 64'h000000000000067F;
assign u[4'b1010] [64] = 64'h0000000000000A7F;
assign v[4'b1010] [64] = 64'h0000000000000E7F;
assign X[4'b1011] [01] = 64'h00000000000002C0;
assign Y[4'b1011] [01] = 64'h0000000000000680;
assign u[4'b1011] [01] = 64'h0000000000000A80;
assign v[4'b1011] [01] = 64'h0000000000000E80;
assign X[4'b1011] [02] = 64'h00000000000002C1;
assign Y[4'b1011] [02] = 64'h0000000000000681;
assign u[4'b1011] [02] = 64'h0000000000000A81;
assign v[4'b1011] [02] = 64'h0000000000000E81;
assign X[4'b1011] [03] = 64'h00000000000002C2;
assign Y[4'b1011] [03] = 64'h0000000000000682;
assign u[4'b1011] [03] = 64'h0000000000000A82;
assign v[4'b1011] [03] = 64'h0000000000000E82;
assign X[4'b1011] [04] = 64'h00000000000002C3;
assign Y[4'b1011] [04] = 64'h0000000000000683;
assign u[4'b1011] [04] = 64'h0000000000000A83;
assign v[4'b1011] [04] = 64'h0000000000000E83;
assign X[4'b1011] [05] = 64'h00000000000002C4;
assign Y[4'b1011] [05] = 64'h0000000000000684;
assign u[4'b1011] [05] = 64'h0000000000000A84;
assign v[4'b1011] [05] = 64'h0000000000000E84;
assign X[4'b1011] [06] = 64'h00000000000002C5;
assign Y[4'b1011] [06] = 64'h0000000000000685;
assign u[4'b1011] [06] = 64'h0000000000000A85;
assign v[4'b1011] [06] = 64'h0000000000000E85;
assign X[4'b1011] [07] = 64'h00000000000002C6;
assign Y[4'b1011] [07] = 64'h0000000000000686;
assign u[4'b1011] [07] = 64'h0000000000000A86;
assign v[4'b1011] [07] = 64'h0000000000000E86;
assign X[4'b1011] [08] = 64'h00000000000002C7;
assign Y[4'b1011] [08] = 64'h0000000000000687;
assign u[4'b1011] [08] = 64'h0000000000000A87;
assign v[4'b1011] [08] = 64'h0000000000000E87;
assign X[4'b1011] [09] = 64'h00000000000002C8;
assign Y[4'b1011] [09] = 64'h0000000000000688;
assign u[4'b1011] [09] = 64'h0000000000000A88;
assign v[4'b1011] [09] = 64'h0000000000000E88;
assign X[4'b1011] [10] = 64'h00000000000002C9;
assign Y[4'b1011] [10] = 64'h0000000000000689;
assign u[4'b1011] [10] = 64'h0000000000000A89;
assign v[4'b1011] [10] = 64'h0000000000000E89;
assign X[4'b1011] [11] = 64'h00000000000002CA;
assign Y[4'b1011] [11] = 64'h000000000000068A;
assign u[4'b1011] [11] = 64'h0000000000000A8A;
assign v[4'b1011] [11] = 64'h0000000000000E8A;
assign X[4'b1011] [12] = 64'h00000000000002CB;
assign Y[4'b1011] [12] = 64'h000000000000068B;
assign u[4'b1011] [12] = 64'h0000000000000A8B;
assign v[4'b1011] [12] = 64'h0000000000000E8B;
assign X[4'b1011] [13] = 64'h00000000000002CC;
assign Y[4'b1011] [13] = 64'h000000000000068C;
assign u[4'b1011] [13] = 64'h0000000000000A8C;
assign v[4'b1011] [13] = 64'h0000000000000E8C;
assign X[4'b1011] [14] = 64'h00000000000002CD;
assign Y[4'b1011] [14] = 64'h000000000000068D;
assign u[4'b1011] [14] = 64'h0000000000000A8D;
assign v[4'b1011] [14] = 64'h0000000000000E8D;
assign X[4'b1011] [15] = 64'h00000000000002CE;
assign Y[4'b1011] [15] = 64'h000000000000068E;
assign u[4'b1011] [15] = 64'h0000000000000A8E;
assign v[4'b1011] [15] = 64'h0000000000000E8E;
assign X[4'b1011] [16] = 64'h00000000000002CF;
assign Y[4'b1011] [16] = 64'h000000000000068F;
assign u[4'b1011] [16] = 64'h0000000000000A8F;
assign v[4'b1011] [16] = 64'h0000000000000E8F;
assign X[4'b1011] [17] = 64'h00000000000002D0;
assign Y[4'b1011] [17] = 64'h0000000000000690;
assign u[4'b1011] [17] = 64'h0000000000000A90;
assign v[4'b1011] [17] = 64'h0000000000000E90;
assign X[4'b1011] [18] = 64'h00000000000002D1;
assign Y[4'b1011] [18] = 64'h0000000000000691;
assign u[4'b1011] [18] = 64'h0000000000000A91;
assign v[4'b1011] [18] = 64'h0000000000000E91;
assign X[4'b1011] [19] = 64'h00000000000002D2;
assign Y[4'b1011] [19] = 64'h0000000000000692;
assign u[4'b1011] [19] = 64'h0000000000000A92;
assign v[4'b1011] [19] = 64'h0000000000000E92;
assign X[4'b1011] [20] = 64'h00000000000002D3;
assign Y[4'b1011] [20] = 64'h0000000000000693;
assign u[4'b1011] [20] = 64'h0000000000000A93;
assign v[4'b1011] [20] = 64'h0000000000000E93;
assign X[4'b1011] [21] = 64'h00000000000002D4;
assign Y[4'b1011] [21] = 64'h0000000000000694;
assign u[4'b1011] [21] = 64'h0000000000000A94;
assign v[4'b1011] [21] = 64'h0000000000000E94;
assign X[4'b1011] [22] = 64'h00000000000002D5;
assign Y[4'b1011] [22] = 64'h0000000000000695;
assign u[4'b1011] [22] = 64'h0000000000000A95;
assign v[4'b1011] [22] = 64'h0000000000000E95;
assign X[4'b1011] [23] = 64'h00000000000002D6;
assign Y[4'b1011] [23] = 64'h0000000000000696;
assign u[4'b1011] [23] = 64'h0000000000000A96;
assign v[4'b1011] [23] = 64'h0000000000000E96;
assign X[4'b1011] [24] = 64'h00000000000002D7;
assign Y[4'b1011] [24] = 64'h0000000000000697;
assign u[4'b1011] [24] = 64'h0000000000000A97;
assign v[4'b1011] [24] = 64'h0000000000000E97;
assign X[4'b1011] [25] = 64'h00000000000002D8;
assign Y[4'b1011] [25] = 64'h0000000000000698;
assign u[4'b1011] [25] = 64'h0000000000000A98;
assign v[4'b1011] [25] = 64'h0000000000000E98;
assign X[4'b1011] [26] = 64'h00000000000002D9;
assign Y[4'b1011] [26] = 64'h0000000000000699;
assign u[4'b1011] [26] = 64'h0000000000000A99;
assign v[4'b1011] [26] = 64'h0000000000000E99;
assign X[4'b1011] [27] = 64'h00000000000002DA;
assign Y[4'b1011] [27] = 64'h000000000000069A;
assign u[4'b1011] [27] = 64'h0000000000000A9A;
assign v[4'b1011] [27] = 64'h0000000000000E9A;
assign X[4'b1011] [28] = 64'h00000000000002DB;
assign Y[4'b1011] [28] = 64'h000000000000069B;
assign u[4'b1011] [28] = 64'h0000000000000A9B;
assign v[4'b1011] [28] = 64'h0000000000000E9B;
assign X[4'b1011] [29] = 64'h00000000000002DC;
assign Y[4'b1011] [29] = 64'h000000000000069C;
assign u[4'b1011] [29] = 64'h0000000000000A9C;
assign v[4'b1011] [29] = 64'h0000000000000E9C;
assign X[4'b1011] [30] = 64'h00000000000002DD;
assign Y[4'b1011] [30] = 64'h000000000000069D;
assign u[4'b1011] [30] = 64'h0000000000000A9D;
assign v[4'b1011] [30] = 64'h0000000000000E9D;
assign X[4'b1011] [31] = 64'h00000000000002DE;
assign Y[4'b1011] [31] = 64'h000000000000069E;
assign u[4'b1011] [31] = 64'h0000000000000A9E;
assign v[4'b1011] [31] = 64'h0000000000000E9E;
assign X[4'b1011] [32] = 64'h00000000000002DF;
assign Y[4'b1011] [32] = 64'h000000000000069F;
assign u[4'b1011] [32] = 64'h0000000000000A9F;
assign v[4'b1011] [32] = 64'h0000000000000E9F;
assign X[4'b1011] [33] = 64'h00000000000002E0;
assign Y[4'b1011] [33] = 64'h00000000000006A0;
assign u[4'b1011] [33] = 64'h0000000000000AA0;
assign v[4'b1011] [33] = 64'h0000000000000EA0;
assign X[4'b1011] [34] = 64'h00000000000002E1;
assign Y[4'b1011] [34] = 64'h00000000000006A1;
assign u[4'b1011] [34] = 64'h0000000000000AA1;
assign v[4'b1011] [34] = 64'h0000000000000EA1;
assign X[4'b1011] [35] = 64'h00000000000002E2;
assign Y[4'b1011] [35] = 64'h00000000000006A2;
assign u[4'b1011] [35] = 64'h0000000000000AA2;
assign v[4'b1011] [35] = 64'h0000000000000EA2;
assign X[4'b1011] [36] = 64'h00000000000002E3;
assign Y[4'b1011] [36] = 64'h00000000000006A3;
assign u[4'b1011] [36] = 64'h0000000000000AA3;
assign v[4'b1011] [36] = 64'h0000000000000EA3;
assign X[4'b1011] [37] = 64'h00000000000002E4;
assign Y[4'b1011] [37] = 64'h00000000000006A4;
assign u[4'b1011] [37] = 64'h0000000000000AA4;
assign v[4'b1011] [37] = 64'h0000000000000EA4;
assign X[4'b1011] [38] = 64'h00000000000002E5;
assign Y[4'b1011] [38] = 64'h00000000000006A5;
assign u[4'b1011] [38] = 64'h0000000000000AA5;
assign v[4'b1011] [38] = 64'h0000000000000EA5;
assign X[4'b1011] [39] = 64'h00000000000002E6;
assign Y[4'b1011] [39] = 64'h00000000000006A6;
assign u[4'b1011] [39] = 64'h0000000000000AA6;
assign v[4'b1011] [39] = 64'h0000000000000EA6;
assign X[4'b1011] [40] = 64'h00000000000002E7;
assign Y[4'b1011] [40] = 64'h00000000000006A7;
assign u[4'b1011] [40] = 64'h0000000000000AA7;
assign v[4'b1011] [40] = 64'h0000000000000EA7;
assign X[4'b1011] [41] = 64'h00000000000002E8;
assign Y[4'b1011] [41] = 64'h00000000000006A8;
assign u[4'b1011] [41] = 64'h0000000000000AA8;
assign v[4'b1011] [41] = 64'h0000000000000EA8;
assign X[4'b1011] [42] = 64'h00000000000002E9;
assign Y[4'b1011] [42] = 64'h00000000000006A9;
assign u[4'b1011] [42] = 64'h0000000000000AA9;
assign v[4'b1011] [42] = 64'h0000000000000EA9;
assign X[4'b1011] [43] = 64'h00000000000002EA;
assign Y[4'b1011] [43] = 64'h00000000000006AA;
assign u[4'b1011] [43] = 64'h0000000000000AAA;
assign v[4'b1011] [43] = 64'h0000000000000EAA;
assign X[4'b1011] [44] = 64'h00000000000002EB;
assign Y[4'b1011] [44] = 64'h00000000000006AB;
assign u[4'b1011] [44] = 64'h0000000000000AAB;
assign v[4'b1011] [44] = 64'h0000000000000EAB;
assign X[4'b1011] [45] = 64'h00000000000002EC;
assign Y[4'b1011] [45] = 64'h00000000000006AC;
assign u[4'b1011] [45] = 64'h0000000000000AAC;
assign v[4'b1011] [45] = 64'h0000000000000EAC;
assign X[4'b1011] [46] = 64'h00000000000002ED;
assign Y[4'b1011] [46] = 64'h00000000000006AD;
assign u[4'b1011] [46] = 64'h0000000000000AAD;
assign v[4'b1011] [46] = 64'h0000000000000EAD;
assign X[4'b1011] [47] = 64'h00000000000002EE;
assign Y[4'b1011] [47] = 64'h00000000000006AE;
assign u[4'b1011] [47] = 64'h0000000000000AAE;
assign v[4'b1011] [47] = 64'h0000000000000EAE;
assign X[4'b1011] [48] = 64'h00000000000002EF;
assign Y[4'b1011] [48] = 64'h00000000000006AF;
assign u[4'b1011] [48] = 64'h0000000000000AAF;
assign v[4'b1011] [48] = 64'h0000000000000EAF;
assign X[4'b1011] [49] = 64'h00000000000002F0;
assign Y[4'b1011] [49] = 64'h00000000000006B0;
assign u[4'b1011] [49] = 64'h0000000000000AB0;
assign v[4'b1011] [49] = 64'h0000000000000EB0;
assign X[4'b1011] [50] = 64'h00000000000002F1;
assign Y[4'b1011] [50] = 64'h00000000000006B1;
assign u[4'b1011] [50] = 64'h0000000000000AB1;
assign v[4'b1011] [50] = 64'h0000000000000EB1;
assign X[4'b1011] [51] = 64'h00000000000002F2;
assign Y[4'b1011] [51] = 64'h00000000000006B2;
assign u[4'b1011] [51] = 64'h0000000000000AB2;
assign v[4'b1011] [51] = 64'h0000000000000EB2;
assign X[4'b1011] [52] = 64'h00000000000002F3;
assign Y[4'b1011] [52] = 64'h00000000000006B3;
assign u[4'b1011] [52] = 64'h0000000000000AB3;
assign v[4'b1011] [52] = 64'h0000000000000EB3;
assign X[4'b1011] [53] = 64'h00000000000002F4;
assign Y[4'b1011] [53] = 64'h00000000000006B4;
assign u[4'b1011] [53] = 64'h0000000000000AB4;
assign v[4'b1011] [53] = 64'h0000000000000EB4;
assign X[4'b1011] [54] = 64'h00000000000002F5;
assign Y[4'b1011] [54] = 64'h00000000000006B5;
assign u[4'b1011] [54] = 64'h0000000000000AB5;
assign v[4'b1011] [54] = 64'h0000000000000EB5;
assign X[4'b1011] [55] = 64'h00000000000002F6;
assign Y[4'b1011] [55] = 64'h00000000000006B6;
assign u[4'b1011] [55] = 64'h0000000000000AB6;
assign v[4'b1011] [55] = 64'h0000000000000EB6;
assign X[4'b1011] [56] = 64'h00000000000002F7;
assign Y[4'b1011] [56] = 64'h00000000000006B7;
assign u[4'b1011] [56] = 64'h0000000000000AB7;
assign v[4'b1011] [56] = 64'h0000000000000EB7;
assign X[4'b1011] [57] = 64'h00000000000002F8;
assign Y[4'b1011] [57] = 64'h00000000000006B8;
assign u[4'b1011] [57] = 64'h0000000000000AB8;
assign v[4'b1011] [57] = 64'h0000000000000EB8;
assign X[4'b1011] [58] = 64'h00000000000002F9;
assign Y[4'b1011] [58] = 64'h00000000000006B9;
assign u[4'b1011] [58] = 64'h0000000000000AB9;
assign v[4'b1011] [58] = 64'h0000000000000EB9;
assign X[4'b1011] [59] = 64'h00000000000002FA;
assign Y[4'b1011] [59] = 64'h00000000000006BA;
assign u[4'b1011] [59] = 64'h0000000000000ABA;
assign v[4'b1011] [59] = 64'h0000000000000EBA;
assign X[4'b1011] [60] = 64'h00000000000002FB;
assign Y[4'b1011] [60] = 64'h00000000000006BB;
assign u[4'b1011] [60] = 64'h0000000000000ABB;
assign v[4'b1011] [60] = 64'h0000000000000EBB;
assign X[4'b1011] [61] = 64'h00000000000002FC;
assign Y[4'b1011] [61] = 64'h00000000000006BC;
assign u[4'b1011] [61] = 64'h0000000000000ABC;
assign v[4'b1011] [61] = 64'h0000000000000EBC;
assign X[4'b1011] [62] = 64'h00000000000002FD;
assign Y[4'b1011] [62] = 64'h00000000000006BD;
assign u[4'b1011] [62] = 64'h0000000000000ABD;
assign v[4'b1011] [62] = 64'h0000000000000EBD;
assign X[4'b1011] [63] = 64'h00000000000002FE;
assign Y[4'b1011] [63] = 64'h00000000000006BE;
assign u[4'b1011] [63] = 64'h0000000000000ABE;
assign v[4'b1011] [63] = 64'h0000000000000EBE;
assign X[4'b1011] [64] = 64'h00000000000002FF;
assign Y[4'b1011] [64] = 64'h00000000000006BF;
assign u[4'b1011] [64] = 64'h0000000000000ABF;
assign v[4'b1011] [64] = 64'h0000000000000EBF;
assign X[4'b1100] [01] = 64'h0000000000000300;
assign Y[4'b1100] [01] = 64'h00000000000006C0;
assign u[4'b1100] [01] = 64'h0000000000000AC0;
assign v[4'b1100] [01] = 64'h0000000000000EC0;
assign X[4'b1100] [02] = 64'h0000000000000301;
assign Y[4'b1100] [02] = 64'h00000000000006C1;
assign u[4'b1100] [02] = 64'h0000000000000AC1;
assign v[4'b1100] [02] = 64'h0000000000000EC1;
assign X[4'b1100] [03] = 64'h0000000000000302;
assign Y[4'b1100] [03] = 64'h00000000000006C2;
assign u[4'b1100] [03] = 64'h0000000000000AC2;
assign v[4'b1100] [03] = 64'h0000000000000EC2;
assign X[4'b1100] [04] = 64'h0000000000000303;
assign Y[4'b1100] [04] = 64'h00000000000006C3;
assign u[4'b1100] [04] = 64'h0000000000000AC3;
assign v[4'b1100] [04] = 64'h0000000000000EC3;
assign X[4'b1100] [05] = 64'h0000000000000304;
assign Y[4'b1100] [05] = 64'h00000000000006C4;
assign u[4'b1100] [05] = 64'h0000000000000AC4;
assign v[4'b1100] [05] = 64'h0000000000000EC4;
assign X[4'b1100] [06] = 64'h0000000000000305;
assign Y[4'b1100] [06] = 64'h00000000000006C5;
assign u[4'b1100] [06] = 64'h0000000000000AC5;
assign v[4'b1100] [06] = 64'h0000000000000EC5;
assign X[4'b1100] [07] = 64'h0000000000000306;
assign Y[4'b1100] [07] = 64'h00000000000006C6;
assign u[4'b1100] [07] = 64'h0000000000000AC6;
assign v[4'b1100] [07] = 64'h0000000000000EC6;
assign X[4'b1100] [08] = 64'h0000000000000307;
assign Y[4'b1100] [08] = 64'h00000000000006C7;
assign u[4'b1100] [08] = 64'h0000000000000AC7;
assign v[4'b1100] [08] = 64'h0000000000000EC7;
assign X[4'b1100] [09] = 64'h0000000000000308;
assign Y[4'b1100] [09] = 64'h00000000000006C8;
assign u[4'b1100] [09] = 64'h0000000000000AC8;
assign v[4'b1100] [09] = 64'h0000000000000EC8;
assign X[4'b1100] [10] = 64'h0000000000000309;
assign Y[4'b1100] [10] = 64'h00000000000006C9;
assign u[4'b1100] [10] = 64'h0000000000000AC9;
assign v[4'b1100] [10] = 64'h0000000000000EC9;
assign X[4'b1100] [11] = 64'h000000000000030A;
assign Y[4'b1100] [11] = 64'h00000000000006CA;
assign u[4'b1100] [11] = 64'h0000000000000ACA;
assign v[4'b1100] [11] = 64'h0000000000000ECA;
assign X[4'b1100] [12] = 64'h000000000000030B;
assign Y[4'b1100] [12] = 64'h00000000000006CB;
assign u[4'b1100] [12] = 64'h0000000000000ACB;
assign v[4'b1100] [12] = 64'h0000000000000ECB;
assign X[4'b1100] [13] = 64'h000000000000030C;
assign Y[4'b1100] [13] = 64'h00000000000006CC;
assign u[4'b1100] [13] = 64'h0000000000000ACC;
assign v[4'b1100] [13] = 64'h0000000000000ECC;
assign X[4'b1100] [14] = 64'h000000000000030D;
assign Y[4'b1100] [14] = 64'h00000000000006CD;
assign u[4'b1100] [14] = 64'h0000000000000ACD;
assign v[4'b1100] [14] = 64'h0000000000000ECD;
assign X[4'b1100] [15] = 64'h000000000000030E;
assign Y[4'b1100] [15] = 64'h00000000000006CE;
assign u[4'b1100] [15] = 64'h0000000000000ACE;
assign v[4'b1100] [15] = 64'h0000000000000ECE;
assign X[4'b1100] [16] = 64'h000000000000030F;
assign Y[4'b1100] [16] = 64'h00000000000006CF;
assign u[4'b1100] [16] = 64'h0000000000000ACF;
assign v[4'b1100] [16] = 64'h0000000000000ECF;
assign X[4'b1100] [17] = 64'h0000000000000310;
assign Y[4'b1100] [17] = 64'h00000000000006D0;
assign u[4'b1100] [17] = 64'h0000000000000AD0;
assign v[4'b1100] [17] = 64'h0000000000000ED0;
assign X[4'b1100] [18] = 64'h0000000000000311;
assign Y[4'b1100] [18] = 64'h00000000000006D1;
assign u[4'b1100] [18] = 64'h0000000000000AD1;
assign v[4'b1100] [18] = 64'h0000000000000ED1;
assign X[4'b1100] [19] = 64'h0000000000000312;
assign Y[4'b1100] [19] = 64'h00000000000006D2;
assign u[4'b1100] [19] = 64'h0000000000000AD2;
assign v[4'b1100] [19] = 64'h0000000000000ED2;
assign X[4'b1100] [20] = 64'h0000000000000313;
assign Y[4'b1100] [20] = 64'h00000000000006D3;
assign u[4'b1100] [20] = 64'h0000000000000AD3;
assign v[4'b1100] [20] = 64'h0000000000000ED3;
assign X[4'b1100] [21] = 64'h0000000000000314;
assign Y[4'b1100] [21] = 64'h00000000000006D4;
assign u[4'b1100] [21] = 64'h0000000000000AD4;
assign v[4'b1100] [21] = 64'h0000000000000ED4;
assign X[4'b1100] [22] = 64'h0000000000000315;
assign Y[4'b1100] [22] = 64'h00000000000006D5;
assign u[4'b1100] [22] = 64'h0000000000000AD5;
assign v[4'b1100] [22] = 64'h0000000000000ED5;
assign X[4'b1100] [23] = 64'h0000000000000316;
assign Y[4'b1100] [23] = 64'h00000000000006D6;
assign u[4'b1100] [23] = 64'h0000000000000AD6;
assign v[4'b1100] [23] = 64'h0000000000000ED6;
assign X[4'b1100] [24] = 64'h0000000000000317;
assign Y[4'b1100] [24] = 64'h00000000000006D7;
assign u[4'b1100] [24] = 64'h0000000000000AD7;
assign v[4'b1100] [24] = 64'h0000000000000ED7;
assign X[4'b1100] [25] = 64'h0000000000000318;
assign Y[4'b1100] [25] = 64'h00000000000006D8;
assign u[4'b1100] [25] = 64'h0000000000000AD8;
assign v[4'b1100] [25] = 64'h0000000000000ED8;
assign X[4'b1100] [26] = 64'h0000000000000319;
assign Y[4'b1100] [26] = 64'h00000000000006D9;
assign u[4'b1100] [26] = 64'h0000000000000AD9;
assign v[4'b1100] [26] = 64'h0000000000000ED9;
assign X[4'b1100] [27] = 64'h000000000000031A;
assign Y[4'b1100] [27] = 64'h00000000000006DA;
assign u[4'b1100] [27] = 64'h0000000000000ADA;
assign v[4'b1100] [27] = 64'h0000000000000EDA;
assign X[4'b1100] [28] = 64'h000000000000031B;
assign Y[4'b1100] [28] = 64'h00000000000006DB;
assign u[4'b1100] [28] = 64'h0000000000000ADB;
assign v[4'b1100] [28] = 64'h0000000000000EDB;
assign X[4'b1100] [29] = 64'h000000000000031C;
assign Y[4'b1100] [29] = 64'h00000000000006DC;
assign u[4'b1100] [29] = 64'h0000000000000ADC;
assign v[4'b1100] [29] = 64'h0000000000000EDC;
assign X[4'b1100] [30] = 64'h000000000000031D;
assign Y[4'b1100] [30] = 64'h00000000000006DD;
assign u[4'b1100] [30] = 64'h0000000000000ADD;
assign v[4'b1100] [30] = 64'h0000000000000EDD;
assign X[4'b1100] [31] = 64'h000000000000031E;
assign Y[4'b1100] [31] = 64'h00000000000006DE;
assign u[4'b1100] [31] = 64'h0000000000000ADE;
assign v[4'b1100] [31] = 64'h0000000000000EDE;
assign X[4'b1100] [32] = 64'h000000000000031F;
assign Y[4'b1100] [32] = 64'h00000000000006DF;
assign u[4'b1100] [32] = 64'h0000000000000ADF;
assign v[4'b1100] [32] = 64'h0000000000000EDF;
assign X[4'b1100] [33] = 64'h0000000000000320;
assign Y[4'b1100] [33] = 64'h00000000000006E0;
assign u[4'b1100] [33] = 64'h0000000000000AE0;
assign v[4'b1100] [33] = 64'h0000000000000EE0;
assign X[4'b1100] [34] = 64'h0000000000000321;
assign Y[4'b1100] [34] = 64'h00000000000006E1;
assign u[4'b1100] [34] = 64'h0000000000000AE1;
assign v[4'b1100] [34] = 64'h0000000000000EE1;
assign X[4'b1100] [35] = 64'h0000000000000322;
assign Y[4'b1100] [35] = 64'h00000000000006E2;
assign u[4'b1100] [35] = 64'h0000000000000AE2;
assign v[4'b1100] [35] = 64'h0000000000000EE2;
assign X[4'b1100] [36] = 64'h0000000000000323;
assign Y[4'b1100] [36] = 64'h00000000000006E3;
assign u[4'b1100] [36] = 64'h0000000000000AE3;
assign v[4'b1100] [36] = 64'h0000000000000EE3;
assign X[4'b1100] [37] = 64'h0000000000000324;
assign Y[4'b1100] [37] = 64'h00000000000006E4;
assign u[4'b1100] [37] = 64'h0000000000000AE4;
assign v[4'b1100] [37] = 64'h0000000000000EE4;
assign X[4'b1100] [38] = 64'h0000000000000325;
assign Y[4'b1100] [38] = 64'h00000000000006E5;
assign u[4'b1100] [38] = 64'h0000000000000AE5;
assign v[4'b1100] [38] = 64'h0000000000000EE5;
assign X[4'b1100] [39] = 64'h0000000000000326;
assign Y[4'b1100] [39] = 64'h00000000000006E6;
assign u[4'b1100] [39] = 64'h0000000000000AE6;
assign v[4'b1100] [39] = 64'h0000000000000EE6;
assign X[4'b1100] [40] = 64'h0000000000000327;
assign Y[4'b1100] [40] = 64'h00000000000006E7;
assign u[4'b1100] [40] = 64'h0000000000000AE7;
assign v[4'b1100] [40] = 64'h0000000000000EE7;
assign X[4'b1100] [41] = 64'h0000000000000328;
assign Y[4'b1100] [41] = 64'h00000000000006E8;
assign u[4'b1100] [41] = 64'h0000000000000AE8;
assign v[4'b1100] [41] = 64'h0000000000000EE8;
assign X[4'b1100] [42] = 64'h0000000000000329;
assign Y[4'b1100] [42] = 64'h00000000000006E9;
assign u[4'b1100] [42] = 64'h0000000000000AE9;
assign v[4'b1100] [42] = 64'h0000000000000EE9;
assign X[4'b1100] [43] = 64'h000000000000032A;
assign Y[4'b1100] [43] = 64'h00000000000006EA;
assign u[4'b1100] [43] = 64'h0000000000000AEA;
assign v[4'b1100] [43] = 64'h0000000000000EEA;
assign X[4'b1100] [44] = 64'h000000000000032B;
assign Y[4'b1100] [44] = 64'h00000000000006EB;
assign u[4'b1100] [44] = 64'h0000000000000AEB;
assign v[4'b1100] [44] = 64'h0000000000000EEB;
assign X[4'b1100] [45] = 64'h000000000000032C;
assign Y[4'b1100] [45] = 64'h00000000000006EC;
assign u[4'b1100] [45] = 64'h0000000000000AEC;
assign v[4'b1100] [45] = 64'h0000000000000EEC;
assign X[4'b1100] [46] = 64'h000000000000032D;
assign Y[4'b1100] [46] = 64'h00000000000006ED;
assign u[4'b1100] [46] = 64'h0000000000000AED;
assign v[4'b1100] [46] = 64'h0000000000000EED;
assign X[4'b1100] [47] = 64'h000000000000032E;
assign Y[4'b1100] [47] = 64'h00000000000006EE;
assign u[4'b1100] [47] = 64'h0000000000000AEE;
assign v[4'b1100] [47] = 64'h0000000000000EEE;
assign X[4'b1100] [48] = 64'h000000000000032F;
assign Y[4'b1100] [48] = 64'h00000000000006EF;
assign u[4'b1100] [48] = 64'h0000000000000AEF;
assign v[4'b1100] [48] = 64'h0000000000000EEF;
assign X[4'b1100] [49] = 64'h0000000000000330;
assign Y[4'b1100] [49] = 64'h00000000000006F0;
assign u[4'b1100] [49] = 64'h0000000000000AF0;
assign v[4'b1100] [49] = 64'h0000000000000EF0;
assign X[4'b1100] [50] = 64'h0000000000000331;
assign Y[4'b1100] [50] = 64'h00000000000006F1;
assign u[4'b1100] [50] = 64'h0000000000000AF1;
assign v[4'b1100] [50] = 64'h0000000000000EF1;
assign X[4'b1100] [51] = 64'h0000000000000332;
assign Y[4'b1100] [51] = 64'h00000000000006F2;
assign u[4'b1100] [51] = 64'h0000000000000AF2;
assign v[4'b1100] [51] = 64'h0000000000000EF2;
assign X[4'b1100] [52] = 64'h0000000000000333;
assign Y[4'b1100] [52] = 64'h00000000000006F3;
assign u[4'b1100] [52] = 64'h0000000000000AF3;
assign v[4'b1100] [52] = 64'h0000000000000EF3;
assign X[4'b1100] [53] = 64'h0000000000000334;
assign Y[4'b1100] [53] = 64'h00000000000006F4;
assign u[4'b1100] [53] = 64'h0000000000000AF4;
assign v[4'b1100] [53] = 64'h0000000000000EF4;
assign X[4'b1100] [54] = 64'h0000000000000335;
assign Y[4'b1100] [54] = 64'h00000000000006F5;
assign u[4'b1100] [54] = 64'h0000000000000AF5;
assign v[4'b1100] [54] = 64'h0000000000000EF5;
assign X[4'b1100] [55] = 64'h0000000000000336;
assign Y[4'b1100] [55] = 64'h00000000000006F6;
assign u[4'b1100] [55] = 64'h0000000000000AF6;
assign v[4'b1100] [55] = 64'h0000000000000EF6;
assign X[4'b1100] [56] = 64'h0000000000000337;
assign Y[4'b1100] [56] = 64'h00000000000006F7;
assign u[4'b1100] [56] = 64'h0000000000000AF7;
assign v[4'b1100] [56] = 64'h0000000000000EF7;
assign X[4'b1100] [57] = 64'h0000000000000338;
assign Y[4'b1100] [57] = 64'h00000000000006F8;
assign u[4'b1100] [57] = 64'h0000000000000AF8;
assign v[4'b1100] [57] = 64'h0000000000000EF8;
assign X[4'b1100] [58] = 64'h0000000000000339;
assign Y[4'b1100] [58] = 64'h00000000000006F9;
assign u[4'b1100] [58] = 64'h0000000000000AF9;
assign v[4'b1100] [58] = 64'h0000000000000EF9;
assign X[4'b1100] [59] = 64'h000000000000033A;
assign Y[4'b1100] [59] = 64'h00000000000006FA;
assign u[4'b1100] [59] = 64'h0000000000000AFA;
assign v[4'b1100] [59] = 64'h0000000000000EFA;
assign X[4'b1100] [60] = 64'h000000000000033B;
assign Y[4'b1100] [60] = 64'h00000000000006FB;
assign u[4'b1100] [60] = 64'h0000000000000AFB;
assign v[4'b1100] [60] = 64'h0000000000000EFB;
assign X[4'b1100] [61] = 64'h000000000000033C;
assign Y[4'b1100] [61] = 64'h00000000000006FC;
assign u[4'b1100] [61] = 64'h0000000000000AFC;
assign v[4'b1100] [61] = 64'h0000000000000EFC;
assign X[4'b1100] [62] = 64'h000000000000033D;
assign Y[4'b1100] [62] = 64'h00000000000006FD;
assign u[4'b1100] [62] = 64'h0000000000000AFD;
assign v[4'b1100] [62] = 64'h0000000000000EFD;
assign X[4'b1100] [63] = 64'h000000000000033E;
assign Y[4'b1100] [63] = 64'h00000000000006FE;
assign u[4'b1100] [63] = 64'h0000000000000AFE;
assign v[4'b1100] [63] = 64'h0000000000000EFE;
assign X[4'b1100] [64] = 64'h000000000000033F;
assign Y[4'b1100] [64] = 64'h00000000000006FF;
assign u[4'b1100] [64] = 64'h0000000000000AFF;
assign v[4'b1100] [64] = 64'h0000000000000EFF;
assign X[4'b1101] [01] = 64'h0000000000000340;
assign Y[4'b1101] [01] = 64'h0000000000000700;
assign u[4'b1101] [01] = 64'h0000000000000B00;
assign v[4'b1101] [01] = 64'h0000000000000F00;
assign X[4'b1101] [02] = 64'h0000000000000341;
assign Y[4'b1101] [02] = 64'h0000000000000701;
assign u[4'b1101] [02] = 64'h0000000000000B01;
assign v[4'b1101] [02] = 64'h0000000000000F01;
assign X[4'b1101] [03] = 64'h0000000000000342;
assign Y[4'b1101] [03] = 64'h0000000000000702;
assign u[4'b1101] [03] = 64'h0000000000000B02;
assign v[4'b1101] [03] = 64'h0000000000000F02;
assign X[4'b1101] [04] = 64'h0000000000000343;
assign Y[4'b1101] [04] = 64'h0000000000000703;
assign u[4'b1101] [04] = 64'h0000000000000B03;
assign v[4'b1101] [04] = 64'h0000000000000F03;
assign X[4'b1101] [05] = 64'h0000000000000344;
assign Y[4'b1101] [05] = 64'h0000000000000704;
assign u[4'b1101] [05] = 64'h0000000000000B04;
assign v[4'b1101] [05] = 64'h0000000000000F04;
assign X[4'b1101] [06] = 64'h0000000000000345;
assign Y[4'b1101] [06] = 64'h0000000000000705;
assign u[4'b1101] [06] = 64'h0000000000000B05;
assign v[4'b1101] [06] = 64'h0000000000000F05;
assign X[4'b1101] [07] = 64'h0000000000000346;
assign Y[4'b1101] [07] = 64'h0000000000000706;
assign u[4'b1101] [07] = 64'h0000000000000B06;
assign v[4'b1101] [07] = 64'h0000000000000F06;
assign X[4'b1101] [08] = 64'h0000000000000347;
assign Y[4'b1101] [08] = 64'h0000000000000707;
assign u[4'b1101] [08] = 64'h0000000000000B07;
assign v[4'b1101] [08] = 64'h0000000000000F07;
assign X[4'b1101] [09] = 64'h0000000000000348;
assign Y[4'b1101] [09] = 64'h0000000000000708;
assign u[4'b1101] [09] = 64'h0000000000000B08;
assign v[4'b1101] [09] = 64'h0000000000000F08;
assign X[4'b1101] [10] = 64'h0000000000000349;
assign Y[4'b1101] [10] = 64'h0000000000000709;
assign u[4'b1101] [10] = 64'h0000000000000B09;
assign v[4'b1101] [10] = 64'h0000000000000F09;
assign X[4'b1101] [11] = 64'h000000000000034A;
assign Y[4'b1101] [11] = 64'h000000000000070A;
assign u[4'b1101] [11] = 64'h0000000000000B0A;
assign v[4'b1101] [11] = 64'h0000000000000F0A;
assign X[4'b1101] [12] = 64'h000000000000034B;
assign Y[4'b1101] [12] = 64'h000000000000070B;
assign u[4'b1101] [12] = 64'h0000000000000B0B;
assign v[4'b1101] [12] = 64'h0000000000000F0B;
assign X[4'b1101] [13] = 64'h000000000000034C;
assign Y[4'b1101] [13] = 64'h000000000000070C;
assign u[4'b1101] [13] = 64'h0000000000000B0C;
assign v[4'b1101] [13] = 64'h0000000000000F0C;
assign X[4'b1101] [14] = 64'h000000000000034D;
assign Y[4'b1101] [14] = 64'h000000000000070D;
assign u[4'b1101] [14] = 64'h0000000000000B0D;
assign v[4'b1101] [14] = 64'h0000000000000F0D;
assign X[4'b1101] [15] = 64'h000000000000034E;
assign Y[4'b1101] [15] = 64'h000000000000070E;
assign u[4'b1101] [15] = 64'h0000000000000B0E;
assign v[4'b1101] [15] = 64'h0000000000000F0E;
assign X[4'b1101] [16] = 64'h000000000000034F;
assign Y[4'b1101] [16] = 64'h000000000000070F;
assign u[4'b1101] [16] = 64'h0000000000000B0F;
assign v[4'b1101] [16] = 64'h0000000000000F0F;
assign X[4'b1101] [17] = 64'h0000000000000350;
assign Y[4'b1101] [17] = 64'h0000000000000710;
assign u[4'b1101] [17] = 64'h0000000000000B10;
assign v[4'b1101] [17] = 64'h0000000000000F10;
assign X[4'b1101] [18] = 64'h0000000000000351;
assign Y[4'b1101] [18] = 64'h0000000000000711;
assign u[4'b1101] [18] = 64'h0000000000000B11;
assign v[4'b1101] [18] = 64'h0000000000000F11;
assign X[4'b1101] [19] = 64'h0000000000000352;
assign Y[4'b1101] [19] = 64'h0000000000000712;
assign u[4'b1101] [19] = 64'h0000000000000B12;
assign v[4'b1101] [19] = 64'h0000000000000F12;
assign X[4'b1101] [20] = 64'h0000000000000353;
assign Y[4'b1101] [20] = 64'h0000000000000713;
assign u[4'b1101] [20] = 64'h0000000000000B13;
assign v[4'b1101] [20] = 64'h0000000000000F13;
assign X[4'b1101] [21] = 64'h0000000000000354;
assign Y[4'b1101] [21] = 64'h0000000000000714;
assign u[4'b1101] [21] = 64'h0000000000000B14;
assign v[4'b1101] [21] = 64'h0000000000000F14;
assign X[4'b1101] [22] = 64'h0000000000000355;
assign Y[4'b1101] [22] = 64'h0000000000000715;
assign u[4'b1101] [22] = 64'h0000000000000B15;
assign v[4'b1101] [22] = 64'h0000000000000F15;
assign X[4'b1101] [23] = 64'h0000000000000356;
assign Y[4'b1101] [23] = 64'h0000000000000716;
assign u[4'b1101] [23] = 64'h0000000000000B16;
assign v[4'b1101] [23] = 64'h0000000000000F16;
assign X[4'b1101] [24] = 64'h0000000000000357;
assign Y[4'b1101] [24] = 64'h0000000000000717;
assign u[4'b1101] [24] = 64'h0000000000000B17;
assign v[4'b1101] [24] = 64'h0000000000000F17;
assign X[4'b1101] [25] = 64'h0000000000000358;
assign Y[4'b1101] [25] = 64'h0000000000000718;
assign u[4'b1101] [25] = 64'h0000000000000B18;
assign v[4'b1101] [25] = 64'h0000000000000F18;
assign X[4'b1101] [26] = 64'h0000000000000359;
assign Y[4'b1101] [26] = 64'h0000000000000719;
assign u[4'b1101] [26] = 64'h0000000000000B19;
assign v[4'b1101] [26] = 64'h0000000000000F19;
assign X[4'b1101] [27] = 64'h000000000000035A;
assign Y[4'b1101] [27] = 64'h000000000000071A;
assign u[4'b1101] [27] = 64'h0000000000000B1A;
assign v[4'b1101] [27] = 64'h0000000000000F1A;
assign X[4'b1101] [28] = 64'h000000000000035B;
assign Y[4'b1101] [28] = 64'h000000000000071B;
assign u[4'b1101] [28] = 64'h0000000000000B1B;
assign v[4'b1101] [28] = 64'h0000000000000F1B;
assign X[4'b1101] [29] = 64'h000000000000035C;
assign Y[4'b1101] [29] = 64'h000000000000071C;
assign u[4'b1101] [29] = 64'h0000000000000B1C;
assign v[4'b1101] [29] = 64'h0000000000000F1C;
assign X[4'b1101] [30] = 64'h000000000000035D;
assign Y[4'b1101] [30] = 64'h000000000000071D;
assign u[4'b1101] [30] = 64'h0000000000000B1D;
assign v[4'b1101] [30] = 64'h0000000000000F1D;
assign X[4'b1101] [31] = 64'h000000000000035E;
assign Y[4'b1101] [31] = 64'h000000000000071E;
assign u[4'b1101] [31] = 64'h0000000000000B1E;
assign v[4'b1101] [31] = 64'h0000000000000F1E;
assign X[4'b1101] [32] = 64'h000000000000035F;
assign Y[4'b1101] [32] = 64'h000000000000071F;
assign u[4'b1101] [32] = 64'h0000000000000B1F;
assign v[4'b1101] [32] = 64'h0000000000000F1F;
assign X[4'b1101] [33] = 64'h0000000000000360;
assign Y[4'b1101] [33] = 64'h0000000000000720;
assign u[4'b1101] [33] = 64'h0000000000000B20;
assign v[4'b1101] [33] = 64'h0000000000000F20;
assign X[4'b1101] [34] = 64'h0000000000000361;
assign Y[4'b1101] [34] = 64'h0000000000000721;
assign u[4'b1101] [34] = 64'h0000000000000B21;
assign v[4'b1101] [34] = 64'h0000000000000F21;
assign X[4'b1101] [35] = 64'h0000000000000362;
assign Y[4'b1101] [35] = 64'h0000000000000722;
assign u[4'b1101] [35] = 64'h0000000000000B22;
assign v[4'b1101] [35] = 64'h0000000000000F22;
assign X[4'b1101] [36] = 64'h0000000000000363;
assign Y[4'b1101] [36] = 64'h0000000000000723;
assign u[4'b1101] [36] = 64'h0000000000000B23;
assign v[4'b1101] [36] = 64'h0000000000000F23;
assign X[4'b1101] [37] = 64'h0000000000000364;
assign Y[4'b1101] [37] = 64'h0000000000000724;
assign u[4'b1101] [37] = 64'h0000000000000B24;
assign v[4'b1101] [37] = 64'h0000000000000F24;
assign X[4'b1101] [38] = 64'h0000000000000365;
assign Y[4'b1101] [38] = 64'h0000000000000725;
assign u[4'b1101] [38] = 64'h0000000000000B25;
assign v[4'b1101] [38] = 64'h0000000000000F25;
assign X[4'b1101] [39] = 64'h0000000000000366;
assign Y[4'b1101] [39] = 64'h0000000000000726;
assign u[4'b1101] [39] = 64'h0000000000000B26;
assign v[4'b1101] [39] = 64'h0000000000000F26;
assign X[4'b1101] [40] = 64'h0000000000000367;
assign Y[4'b1101] [40] = 64'h0000000000000727;
assign u[4'b1101] [40] = 64'h0000000000000B27;
assign v[4'b1101] [40] = 64'h0000000000000F27;
assign X[4'b1101] [41] = 64'h0000000000000368;
assign Y[4'b1101] [41] = 64'h0000000000000728;
assign u[4'b1101] [41] = 64'h0000000000000B28;
assign v[4'b1101] [41] = 64'h0000000000000F28;
assign X[4'b1101] [42] = 64'h0000000000000369;
assign Y[4'b1101] [42] = 64'h0000000000000729;
assign u[4'b1101] [42] = 64'h0000000000000B29;
assign v[4'b1101] [42] = 64'h0000000000000F29;
assign X[4'b1101] [43] = 64'h000000000000036A;
assign Y[4'b1101] [43] = 64'h000000000000072A;
assign u[4'b1101] [43] = 64'h0000000000000B2A;
assign v[4'b1101] [43] = 64'h0000000000000F2A;
assign X[4'b1101] [44] = 64'h000000000000036B;
assign Y[4'b1101] [44] = 64'h000000000000072B;
assign u[4'b1101] [44] = 64'h0000000000000B2B;
assign v[4'b1101] [44] = 64'h0000000000000F2B;
assign X[4'b1101] [45] = 64'h000000000000036C;
assign Y[4'b1101] [45] = 64'h000000000000072C;
assign u[4'b1101] [45] = 64'h0000000000000B2C;
assign v[4'b1101] [45] = 64'h0000000000000F2C;
assign X[4'b1101] [46] = 64'h000000000000036D;
assign Y[4'b1101] [46] = 64'h000000000000072D;
assign u[4'b1101] [46] = 64'h0000000000000B2D;
assign v[4'b1101] [46] = 64'h0000000000000F2D;
assign X[4'b1101] [47] = 64'h000000000000036E;
assign Y[4'b1101] [47] = 64'h000000000000072E;
assign u[4'b1101] [47] = 64'h0000000000000B2E;
assign v[4'b1101] [47] = 64'h0000000000000F2E;
assign X[4'b1101] [48] = 64'h000000000000036F;
assign Y[4'b1101] [48] = 64'h000000000000072F;
assign u[4'b1101] [48] = 64'h0000000000000B2F;
assign v[4'b1101] [48] = 64'h0000000000000F2F;
assign X[4'b1101] [49] = 64'h0000000000000370;
assign Y[4'b1101] [49] = 64'h0000000000000730;
assign u[4'b1101] [49] = 64'h0000000000000B30;
assign v[4'b1101] [49] = 64'h0000000000000F30;
assign X[4'b1101] [50] = 64'h0000000000000371;
assign Y[4'b1101] [50] = 64'h0000000000000731;
assign u[4'b1101] [50] = 64'h0000000000000B31;
assign v[4'b1101] [50] = 64'h0000000000000F31;
assign X[4'b1101] [51] = 64'h0000000000000372;
assign Y[4'b1101] [51] = 64'h0000000000000732;
assign u[4'b1101] [51] = 64'h0000000000000B32;
assign v[4'b1101] [51] = 64'h0000000000000F32;
assign X[4'b1101] [52] = 64'h0000000000000373;
assign Y[4'b1101] [52] = 64'h0000000000000733;
assign u[4'b1101] [52] = 64'h0000000000000B33;
assign v[4'b1101] [52] = 64'h0000000000000F33;
assign X[4'b1101] [53] = 64'h0000000000000374;
assign Y[4'b1101] [53] = 64'h0000000000000734;
assign u[4'b1101] [53] = 64'h0000000000000B34;
assign v[4'b1101] [53] = 64'h0000000000000F34;
assign X[4'b1101] [54] = 64'h0000000000000375;
assign Y[4'b1101] [54] = 64'h0000000000000735;
assign u[4'b1101] [54] = 64'h0000000000000B35;
assign v[4'b1101] [54] = 64'h0000000000000F35;
assign X[4'b1101] [55] = 64'h0000000000000376;
assign Y[4'b1101] [55] = 64'h0000000000000736;
assign u[4'b1101] [55] = 64'h0000000000000B36;
assign v[4'b1101] [55] = 64'h0000000000000F36;
assign X[4'b1101] [56] = 64'h0000000000000377;
assign Y[4'b1101] [56] = 64'h0000000000000737;
assign u[4'b1101] [56] = 64'h0000000000000B37;
assign v[4'b1101] [56] = 64'h0000000000000F37;
assign X[4'b1101] [57] = 64'h0000000000000378;
assign Y[4'b1101] [57] = 64'h0000000000000738;
assign u[4'b1101] [57] = 64'h0000000000000B38;
assign v[4'b1101] [57] = 64'h0000000000000F38;
assign X[4'b1101] [58] = 64'h0000000000000379;
assign Y[4'b1101] [58] = 64'h0000000000000739;
assign u[4'b1101] [58] = 64'h0000000000000B39;
assign v[4'b1101] [58] = 64'h0000000000000F39;
assign X[4'b1101] [59] = 64'h000000000000037A;
assign Y[4'b1101] [59] = 64'h000000000000073A;
assign u[4'b1101] [59] = 64'h0000000000000B3A;
assign v[4'b1101] [59] = 64'h0000000000000F3A;
assign X[4'b1101] [60] = 64'h000000000000037B;
assign Y[4'b1101] [60] = 64'h000000000000073B;
assign u[4'b1101] [60] = 64'h0000000000000B3B;
assign v[4'b1101] [60] = 64'h0000000000000F3B;
assign X[4'b1101] [61] = 64'h000000000000037C;
assign Y[4'b1101] [61] = 64'h000000000000073C;
assign u[4'b1101] [61] = 64'h0000000000000B3C;
assign v[4'b1101] [61] = 64'h0000000000000F3C;
assign X[4'b1101] [62] = 64'h000000000000037D;
assign Y[4'b1101] [62] = 64'h000000000000073D;
assign u[4'b1101] [62] = 64'h0000000000000B3D;
assign v[4'b1101] [62] = 64'h0000000000000F3D;
assign X[4'b1101] [63] = 64'h000000000000037E;
assign Y[4'b1101] [63] = 64'h000000000000073E;
assign u[4'b1101] [63] = 64'h0000000000000B3E;
assign v[4'b1101] [63] = 64'h0000000000000F3E;
assign X[4'b1101] [64] = 64'h000000000000037F;
assign Y[4'b1101] [64] = 64'h000000000000073F;
assign u[4'b1101] [64] = 64'h0000000000000B3F;
assign v[4'b1101] [64] = 64'h0000000000000F3F;
assign X[4'b1110] [01] = 64'h0000000000000380;
assign Y[4'b1110] [01] = 64'h0000000000000740;
assign u[4'b1110] [01] = 64'h0000000000000B40;
assign v[4'b1110] [01] = 64'h0000000000000F40;
assign X[4'b1110] [02] = 64'h0000000000000381;
assign Y[4'b1110] [02] = 64'h0000000000000741;
assign u[4'b1110] [02] = 64'h0000000000000B41;
assign v[4'b1110] [02] = 64'h0000000000000F41;
assign X[4'b1110] [03] = 64'h0000000000000382;
assign Y[4'b1110] [03] = 64'h0000000000000742;
assign u[4'b1110] [03] = 64'h0000000000000B42;
assign v[4'b1110] [03] = 64'h0000000000000F42;
assign X[4'b1110] [04] = 64'h0000000000000383;
assign Y[4'b1110] [04] = 64'h0000000000000743;
assign u[4'b1110] [04] = 64'h0000000000000B43;
assign v[4'b1110] [04] = 64'h0000000000000F43;
assign X[4'b1110] [05] = 64'h0000000000000384;
assign Y[4'b1110] [05] = 64'h0000000000000744;
assign u[4'b1110] [05] = 64'h0000000000000B44;
assign v[4'b1110] [05] = 64'h0000000000000F44;
assign X[4'b1110] [06] = 64'h0000000000000385;
assign Y[4'b1110] [06] = 64'h0000000000000745;
assign u[4'b1110] [06] = 64'h0000000000000B45;
assign v[4'b1110] [06] = 64'h0000000000000F45;
assign X[4'b1110] [07] = 64'h0000000000000386;
assign Y[4'b1110] [07] = 64'h0000000000000746;
assign u[4'b1110] [07] = 64'h0000000000000B46;
assign v[4'b1110] [07] = 64'h0000000000000F46;
assign X[4'b1110] [08] = 64'h0000000000000387;
assign Y[4'b1110] [08] = 64'h0000000000000747;
assign u[4'b1110] [08] = 64'h0000000000000B47;
assign v[4'b1110] [08] = 64'h0000000000000F47;
assign X[4'b1110] [09] = 64'h0000000000000388;
assign Y[4'b1110] [09] = 64'h0000000000000748;
assign u[4'b1110] [09] = 64'h0000000000000B48;
assign v[4'b1110] [09] = 64'h0000000000000F48;
assign X[4'b1110] [10] = 64'h0000000000000389;
assign Y[4'b1110] [10] = 64'h0000000000000749;
assign u[4'b1110] [10] = 64'h0000000000000B49;
assign v[4'b1110] [10] = 64'h0000000000000F49;
assign X[4'b1110] [11] = 64'h000000000000038A;
assign Y[4'b1110] [11] = 64'h000000000000074A;
assign u[4'b1110] [11] = 64'h0000000000000B4A;
assign v[4'b1110] [11] = 64'h0000000000000F4A;
assign X[4'b1110] [12] = 64'h000000000000038B;
assign Y[4'b1110] [12] = 64'h000000000000074B;
assign u[4'b1110] [12] = 64'h0000000000000B4B;
assign v[4'b1110] [12] = 64'h0000000000000F4B;
assign X[4'b1110] [13] = 64'h000000000000038C;
assign Y[4'b1110] [13] = 64'h000000000000074C;
assign u[4'b1110] [13] = 64'h0000000000000B4C;
assign v[4'b1110] [13] = 64'h0000000000000F4C;
assign X[4'b1110] [14] = 64'h000000000000038D;
assign Y[4'b1110] [14] = 64'h000000000000074D;
assign u[4'b1110] [14] = 64'h0000000000000B4D;
assign v[4'b1110] [14] = 64'h0000000000000F4D;
assign X[4'b1110] [15] = 64'h000000000000038E;
assign Y[4'b1110] [15] = 64'h000000000000074E;
assign u[4'b1110] [15] = 64'h0000000000000B4E;
assign v[4'b1110] [15] = 64'h0000000000000F4E;
assign X[4'b1110] [16] = 64'h000000000000038F;
assign Y[4'b1110] [16] = 64'h000000000000074F;
assign u[4'b1110] [16] = 64'h0000000000000B4F;
assign v[4'b1110] [16] = 64'h0000000000000F4F;
assign X[4'b1110] [17] = 64'h0000000000000390;
assign Y[4'b1110] [17] = 64'h0000000000000750;
assign u[4'b1110] [17] = 64'h0000000000000B50;
assign v[4'b1110] [17] = 64'h0000000000000F50;
assign X[4'b1110] [18] = 64'h0000000000000391;
assign Y[4'b1110] [18] = 64'h0000000000000751;
assign u[4'b1110] [18] = 64'h0000000000000B51;
assign v[4'b1110] [18] = 64'h0000000000000F51;
assign X[4'b1110] [19] = 64'h0000000000000392;
assign Y[4'b1110] [19] = 64'h0000000000000752;
assign u[4'b1110] [19] = 64'h0000000000000B52;
assign v[4'b1110] [19] = 64'h0000000000000F52;
assign X[4'b1110] [20] = 64'h0000000000000393;
assign Y[4'b1110] [20] = 64'h0000000000000753;
assign u[4'b1110] [20] = 64'h0000000000000B53;
assign v[4'b1110] [20] = 64'h0000000000000F53;
assign X[4'b1110] [21] = 64'h0000000000000394;
assign Y[4'b1110] [21] = 64'h0000000000000754;
assign u[4'b1110] [21] = 64'h0000000000000B54;
assign v[4'b1110] [21] = 64'h0000000000000F54;
assign X[4'b1110] [22] = 64'h0000000000000395;
assign Y[4'b1110] [22] = 64'h0000000000000755;
assign u[4'b1110] [22] = 64'h0000000000000B55;
assign v[4'b1110] [22] = 64'h0000000000000F55;
assign X[4'b1110] [23] = 64'h0000000000000396;
assign Y[4'b1110] [23] = 64'h0000000000000756;
assign u[4'b1110] [23] = 64'h0000000000000B56;
assign v[4'b1110] [23] = 64'h0000000000000F56;
assign X[4'b1110] [24] = 64'h0000000000000397;
assign Y[4'b1110] [24] = 64'h0000000000000757;
assign u[4'b1110] [24] = 64'h0000000000000B57;
assign v[4'b1110] [24] = 64'h0000000000000F57;
assign X[4'b1110] [25] = 64'h0000000000000398;
assign Y[4'b1110] [25] = 64'h0000000000000758;
assign u[4'b1110] [25] = 64'h0000000000000B58;
assign v[4'b1110] [25] = 64'h0000000000000F58;
assign X[4'b1110] [26] = 64'h0000000000000399;
assign Y[4'b1110] [26] = 64'h0000000000000759;
assign u[4'b1110] [26] = 64'h0000000000000B59;
assign v[4'b1110] [26] = 64'h0000000000000F59;
assign X[4'b1110] [27] = 64'h000000000000039A;
assign Y[4'b1110] [27] = 64'h000000000000075A;
assign u[4'b1110] [27] = 64'h0000000000000B5A;
assign v[4'b1110] [27] = 64'h0000000000000F5A;
assign X[4'b1110] [28] = 64'h000000000000039B;
assign Y[4'b1110] [28] = 64'h000000000000075B;
assign u[4'b1110] [28] = 64'h0000000000000B5B;
assign v[4'b1110] [28] = 64'h0000000000000F5B;
assign X[4'b1110] [29] = 64'h000000000000039C;
assign Y[4'b1110] [29] = 64'h000000000000075C;
assign u[4'b1110] [29] = 64'h0000000000000B5C;
assign v[4'b1110] [29] = 64'h0000000000000F5C;
assign X[4'b1110] [30] = 64'h000000000000039D;
assign Y[4'b1110] [30] = 64'h000000000000075D;
assign u[4'b1110] [30] = 64'h0000000000000B5D;
assign v[4'b1110] [30] = 64'h0000000000000F5D;
assign X[4'b1110] [31] = 64'h000000000000039E;
assign Y[4'b1110] [31] = 64'h000000000000075E;
assign u[4'b1110] [31] = 64'h0000000000000B5E;
assign v[4'b1110] [31] = 64'h0000000000000F5E;
assign X[4'b1110] [32] = 64'h000000000000039F;
assign Y[4'b1110] [32] = 64'h000000000000075F;
assign u[4'b1110] [32] = 64'h0000000000000B5F;
assign v[4'b1110] [32] = 64'h0000000000000F5F;
assign X[4'b1110] [33] = 64'h00000000000003A0;
assign Y[4'b1110] [33] = 64'h0000000000000760;
assign u[4'b1110] [33] = 64'h0000000000000B60;
assign v[4'b1110] [33] = 64'h0000000000000F60;
assign X[4'b1110] [34] = 64'h00000000000003A1;
assign Y[4'b1110] [34] = 64'h0000000000000761;
assign u[4'b1110] [34] = 64'h0000000000000B61;
assign v[4'b1110] [34] = 64'h0000000000000F61;
assign X[4'b1110] [35] = 64'h00000000000003A2;
assign Y[4'b1110] [35] = 64'h0000000000000762;
assign u[4'b1110] [35] = 64'h0000000000000B62;
assign v[4'b1110] [35] = 64'h0000000000000F62;
assign X[4'b1110] [36] = 64'h00000000000003A3;
assign Y[4'b1110] [36] = 64'h0000000000000763;
assign u[4'b1110] [36] = 64'h0000000000000B63;
assign v[4'b1110] [36] = 64'h0000000000000F63;
assign X[4'b1110] [37] = 64'h00000000000003A4;
assign Y[4'b1110] [37] = 64'h0000000000000764;
assign u[4'b1110] [37] = 64'h0000000000000B64;
assign v[4'b1110] [37] = 64'h0000000000000F64;
assign X[4'b1110] [38] = 64'h00000000000003A5;
assign Y[4'b1110] [38] = 64'h0000000000000765;
assign u[4'b1110] [38] = 64'h0000000000000B65;
assign v[4'b1110] [38] = 64'h0000000000000F65;
assign X[4'b1110] [39] = 64'h00000000000003A6;
assign Y[4'b1110] [39] = 64'h0000000000000766;
assign u[4'b1110] [39] = 64'h0000000000000B66;
assign v[4'b1110] [39] = 64'h0000000000000F66;
assign X[4'b1110] [40] = 64'h00000000000003A7;
assign Y[4'b1110] [40] = 64'h0000000000000767;
assign u[4'b1110] [40] = 64'h0000000000000B67;
assign v[4'b1110] [40] = 64'h0000000000000F67;
assign X[4'b1110] [41] = 64'h00000000000003A8;
assign Y[4'b1110] [41] = 64'h0000000000000768;
assign u[4'b1110] [41] = 64'h0000000000000B68;
assign v[4'b1110] [41] = 64'h0000000000000F68;
assign X[4'b1110] [42] = 64'h00000000000003A9;
assign Y[4'b1110] [42] = 64'h0000000000000769;
assign u[4'b1110] [42] = 64'h0000000000000B69;
assign v[4'b1110] [42] = 64'h0000000000000F69;
assign X[4'b1110] [43] = 64'h00000000000003AA;
assign Y[4'b1110] [43] = 64'h000000000000076A;
assign u[4'b1110] [43] = 64'h0000000000000B6A;
assign v[4'b1110] [43] = 64'h0000000000000F6A;
assign X[4'b1110] [44] = 64'h00000000000003AB;
assign Y[4'b1110] [44] = 64'h000000000000076B;
assign u[4'b1110] [44] = 64'h0000000000000B6B;
assign v[4'b1110] [44] = 64'h0000000000000F6B;
assign X[4'b1110] [45] = 64'h00000000000003AC;
assign Y[4'b1110] [45] = 64'h000000000000076C;
assign u[4'b1110] [45] = 64'h0000000000000B6C;
assign v[4'b1110] [45] = 64'h0000000000000F6C;
assign X[4'b1110] [46] = 64'h00000000000003AD;
assign Y[4'b1110] [46] = 64'h000000000000076D;
assign u[4'b1110] [46] = 64'h0000000000000B6D;
assign v[4'b1110] [46] = 64'h0000000000000F6D;
assign X[4'b1110] [47] = 64'h00000000000003AE;
assign Y[4'b1110] [47] = 64'h000000000000076E;
assign u[4'b1110] [47] = 64'h0000000000000B6E;
assign v[4'b1110] [47] = 64'h0000000000000F6E;
assign X[4'b1110] [48] = 64'h00000000000003AF;
assign Y[4'b1110] [48] = 64'h000000000000076F;
assign u[4'b1110] [48] = 64'h0000000000000B6F;
assign v[4'b1110] [48] = 64'h0000000000000F6F;
assign X[4'b1110] [49] = 64'h00000000000003B0;
assign Y[4'b1110] [49] = 64'h0000000000000770;
assign u[4'b1110] [49] = 64'h0000000000000B70;
assign v[4'b1110] [49] = 64'h0000000000000F70;
assign X[4'b1110] [50] = 64'h00000000000003B1;
assign Y[4'b1110] [50] = 64'h0000000000000771;
assign u[4'b1110] [50] = 64'h0000000000000B71;
assign v[4'b1110] [50] = 64'h0000000000000F71;
assign X[4'b1110] [51] = 64'h00000000000003B2;
assign Y[4'b1110] [51] = 64'h0000000000000772;
assign u[4'b1110] [51] = 64'h0000000000000B72;
assign v[4'b1110] [51] = 64'h0000000000000F72;
assign X[4'b1110] [52] = 64'h00000000000003B3;
assign Y[4'b1110] [52] = 64'h0000000000000773;
assign u[4'b1110] [52] = 64'h0000000000000B73;
assign v[4'b1110] [52] = 64'h0000000000000F73;
assign X[4'b1110] [53] = 64'h00000000000003B4;
assign Y[4'b1110] [53] = 64'h0000000000000774;
assign u[4'b1110] [53] = 64'h0000000000000B74;
assign v[4'b1110] [53] = 64'h0000000000000F74;
assign X[4'b1110] [54] = 64'h00000000000003B5;
assign Y[4'b1110] [54] = 64'h0000000000000775;
assign u[4'b1110] [54] = 64'h0000000000000B75;
assign v[4'b1110] [54] = 64'h0000000000000F75;
assign X[4'b1110] [55] = 64'h00000000000003B6;
assign Y[4'b1110] [55] = 64'h0000000000000776;
assign u[4'b1110] [55] = 64'h0000000000000B76;
assign v[4'b1110] [55] = 64'h0000000000000F76;
assign X[4'b1110] [56] = 64'h00000000000003B7;
assign Y[4'b1110] [56] = 64'h0000000000000777;
assign u[4'b1110] [56] = 64'h0000000000000B77;
assign v[4'b1110] [56] = 64'h0000000000000F77;
assign X[4'b1110] [57] = 64'h00000000000003B8;
assign Y[4'b1110] [57] = 64'h0000000000000778;
assign u[4'b1110] [57] = 64'h0000000000000B78;
assign v[4'b1110] [57] = 64'h0000000000000F78;
assign X[4'b1110] [58] = 64'h00000000000003B9;
assign Y[4'b1110] [58] = 64'h0000000000000779;
assign u[4'b1110] [58] = 64'h0000000000000B79;
assign v[4'b1110] [58] = 64'h0000000000000F79;
assign X[4'b1110] [59] = 64'h00000000000003BA;
assign Y[4'b1110] [59] = 64'h000000000000077A;
assign u[4'b1110] [59] = 64'h0000000000000B7A;
assign v[4'b1110] [59] = 64'h0000000000000F7A;
assign X[4'b1110] [60] = 64'h00000000000003BB;
assign Y[4'b1110] [60] = 64'h000000000000077B;
assign u[4'b1110] [60] = 64'h0000000000000B7B;
assign v[4'b1110] [60] = 64'h0000000000000F7B;
assign X[4'b1110] [61] = 64'h00000000000003BC;
assign Y[4'b1110] [61] = 64'h000000000000077C;
assign u[4'b1110] [61] = 64'h0000000000000B7C;
assign v[4'b1110] [61] = 64'h0000000000000F7C;
assign X[4'b1110] [62] = 64'h00000000000003BD;
assign Y[4'b1110] [62] = 64'h000000000000077D;
assign u[4'b1110] [62] = 64'h0000000000000B7D;
assign v[4'b1110] [62] = 64'h0000000000000F7D;
assign X[4'b1110] [63] = 64'h00000000000003BE;
assign Y[4'b1110] [63] = 64'h000000000000077E;
assign u[4'b1110] [63] = 64'h0000000000000B7E;
assign v[4'b1110] [63] = 64'h0000000000000F7E;
assign X[4'b1110] [64] = 64'h00000000000003BF;
assign Y[4'b1110] [64] = 64'h000000000000077F;
assign u[4'b1110] [64] = 64'h0000000000000B7F;
assign v[4'b1110] [64] = 64'h0000000000000F7F;
assign X[4'b1111] [01] = 64'h00000000000003C0;
assign Y[4'b1111] [01] = 64'h0000000000000780;
assign u[4'b1111] [01] = 64'h0000000000000B80;
assign v[4'b1111] [01] = 64'h0000000000000F80;
assign X[4'b1111] [02] = 64'h00000000000003C1;
assign Y[4'b1111] [02] = 64'h0000000000000781;
assign u[4'b1111] [02] = 64'h0000000000000B81;
assign v[4'b1111] [02] = 64'h0000000000000F81;
assign X[4'b1111] [03] = 64'h00000000000003C2;
assign Y[4'b1111] [03] = 64'h0000000000000782;
assign u[4'b1111] [03] = 64'h0000000000000B82;
assign v[4'b1111] [03] = 64'h0000000000000F82;
assign X[4'b1111] [04] = 64'h00000000000003C3;
assign Y[4'b1111] [04] = 64'h0000000000000783;
assign u[4'b1111] [04] = 64'h0000000000000B83;
assign v[4'b1111] [04] = 64'h0000000000000F83;
assign X[4'b1111] [05] = 64'h00000000000003C4;
assign Y[4'b1111] [05] = 64'h0000000000000784;
assign u[4'b1111] [05] = 64'h0000000000000B84;
assign v[4'b1111] [05] = 64'h0000000000000F84;
assign X[4'b1111] [06] = 64'h00000000000003C5;
assign Y[4'b1111] [06] = 64'h0000000000000785;
assign u[4'b1111] [06] = 64'h0000000000000B85;
assign v[4'b1111] [06] = 64'h0000000000000F85;
assign X[4'b1111] [07] = 64'h00000000000003C6;
assign Y[4'b1111] [07] = 64'h0000000000000786;
assign u[4'b1111] [07] = 64'h0000000000000B86;
assign v[4'b1111] [07] = 64'h0000000000000F86;
assign X[4'b1111] [08] = 64'h00000000000003C7;
assign Y[4'b1111] [08] = 64'h0000000000000787;
assign u[4'b1111] [08] = 64'h0000000000000B87;
assign v[4'b1111] [08] = 64'h0000000000000F87;
assign X[4'b1111] [09] = 64'h00000000000003C8;
assign Y[4'b1111] [09] = 64'h0000000000000788;
assign u[4'b1111] [09] = 64'h0000000000000B88;
assign v[4'b1111] [09] = 64'h0000000000000F88;
assign X[4'b1111] [10] = 64'h00000000000003C9;
assign Y[4'b1111] [10] = 64'h0000000000000789;
assign u[4'b1111] [10] = 64'h0000000000000B89;
assign v[4'b1111] [10] = 64'h0000000000000F89;
assign X[4'b1111] [11] = 64'h00000000000003CA;
assign Y[4'b1111] [11] = 64'h000000000000078A;
assign u[4'b1111] [11] = 64'h0000000000000B8A;
assign v[4'b1111] [11] = 64'h0000000000000F8A;
assign X[4'b1111] [12] = 64'h00000000000003CB;
assign Y[4'b1111] [12] = 64'h000000000000078B;
assign u[4'b1111] [12] = 64'h0000000000000B8B;
assign v[4'b1111] [12] = 64'h0000000000000F8B;
assign X[4'b1111] [13] = 64'h00000000000003CC;
assign Y[4'b1111] [13] = 64'h000000000000078C;
assign u[4'b1111] [13] = 64'h0000000000000B8C;
assign v[4'b1111] [13] = 64'h0000000000000F8C;
assign X[4'b1111] [14] = 64'h00000000000003CD;
assign Y[4'b1111] [14] = 64'h000000000000078D;
assign u[4'b1111] [14] = 64'h0000000000000B8D;
assign v[4'b1111] [14] = 64'h0000000000000F8D;
assign X[4'b1111] [15] = 64'h00000000000003CE;
assign Y[4'b1111] [15] = 64'h000000000000078E;
assign u[4'b1111] [15] = 64'h0000000000000B8E;
assign v[4'b1111] [15] = 64'h0000000000000F8E;
assign X[4'b1111] [16] = 64'h00000000000003CF;
assign Y[4'b1111] [16] = 64'h000000000000078F;
assign u[4'b1111] [16] = 64'h0000000000000B8F;
assign v[4'b1111] [16] = 64'h0000000000000F8F;
assign X[4'b1111] [17] = 64'h00000000000003D0;
assign Y[4'b1111] [17] = 64'h0000000000000790;
assign u[4'b1111] [17] = 64'h0000000000000B90;
assign v[4'b1111] [17] = 64'h0000000000000F90;
assign X[4'b1111] [18] = 64'h00000000000003D1;
assign Y[4'b1111] [18] = 64'h0000000000000791;
assign u[4'b1111] [18] = 64'h0000000000000B91;
assign v[4'b1111] [18] = 64'h0000000000000F91;
assign X[4'b1111] [19] = 64'h00000000000003D2;
assign Y[4'b1111] [19] = 64'h0000000000000792;
assign u[4'b1111] [19] = 64'h0000000000000B92;
assign v[4'b1111] [19] = 64'h0000000000000F92;
assign X[4'b1111] [20] = 64'h00000000000003D3;
assign Y[4'b1111] [20] = 64'h0000000000000793;
assign u[4'b1111] [20] = 64'h0000000000000B93;
assign v[4'b1111] [20] = 64'h0000000000000F93;
assign X[4'b1111] [21] = 64'h00000000000003D4;
assign Y[4'b1111] [21] = 64'h0000000000000794;
assign u[4'b1111] [21] = 64'h0000000000000B94;
assign v[4'b1111] [21] = 64'h0000000000000F94;
assign X[4'b1111] [22] = 64'h00000000000003D5;
assign Y[4'b1111] [22] = 64'h0000000000000795;
assign u[4'b1111] [22] = 64'h0000000000000B95;
assign v[4'b1111] [22] = 64'h0000000000000F95;
assign X[4'b1111] [23] = 64'h00000000000003D6;
assign Y[4'b1111] [23] = 64'h0000000000000796;
assign u[4'b1111] [23] = 64'h0000000000000B96;
assign v[4'b1111] [23] = 64'h0000000000000F96;
assign X[4'b1111] [24] = 64'h00000000000003D7;
assign Y[4'b1111] [24] = 64'h0000000000000797;
assign u[4'b1111] [24] = 64'h0000000000000B97;
assign v[4'b1111] [24] = 64'h0000000000000F97;
assign X[4'b1111] [25] = 64'h00000000000003D8;
assign Y[4'b1111] [25] = 64'h0000000000000798;
assign u[4'b1111] [25] = 64'h0000000000000B98;
assign v[4'b1111] [25] = 64'h0000000000000F98;
assign X[4'b1111] [26] = 64'h00000000000003D9;
assign Y[4'b1111] [26] = 64'h0000000000000799;
assign u[4'b1111] [26] = 64'h0000000000000B99;
assign v[4'b1111] [26] = 64'h0000000000000F99;
assign X[4'b1111] [27] = 64'h00000000000003DA;
assign Y[4'b1111] [27] = 64'h000000000000079A;
assign u[4'b1111] [27] = 64'h0000000000000B9A;
assign v[4'b1111] [27] = 64'h0000000000000F9A;
assign X[4'b1111] [28] = 64'h00000000000003DB;
assign Y[4'b1111] [28] = 64'h000000000000079B;
assign u[4'b1111] [28] = 64'h0000000000000B9B;
assign v[4'b1111] [28] = 64'h0000000000000F9B;
assign X[4'b1111] [29] = 64'h00000000000003DC;
assign Y[4'b1111] [29] = 64'h000000000000079C;
assign u[4'b1111] [29] = 64'h0000000000000B9C;
assign v[4'b1111] [29] = 64'h0000000000000F9C;
assign X[4'b1111] [30] = 64'h00000000000003DD;
assign Y[4'b1111] [30] = 64'h000000000000079D;
assign u[4'b1111] [30] = 64'h0000000000000B9D;
assign v[4'b1111] [30] = 64'h0000000000000F9D;
assign X[4'b1111] [31] = 64'h00000000000003DE;
assign Y[4'b1111] [31] = 64'h000000000000079E;
assign u[4'b1111] [31] = 64'h0000000000000B9E;
assign v[4'b1111] [31] = 64'h0000000000000F9E;
assign X[4'b1111] [32] = 64'h00000000000003DF;
assign Y[4'b1111] [32] = 64'h000000000000079F;
assign u[4'b1111] [32] = 64'h0000000000000B9F;
assign v[4'b1111] [32] = 64'h0000000000000F9F;
assign X[4'b1111] [33] = 64'h00000000000003E0;
assign Y[4'b1111] [33] = 64'h00000000000007A0;
assign u[4'b1111] [33] = 64'h0000000000000BA0;
assign v[4'b1111] [33] = 64'h0000000000000FA0;
assign X[4'b1111] [34] = 64'h00000000000003E1;
assign Y[4'b1111] [34] = 64'h00000000000007A1;
assign u[4'b1111] [34] = 64'h0000000000000BA1;
assign v[4'b1111] [34] = 64'h0000000000000FA1;
assign X[4'b1111] [35] = 64'h00000000000003E2;
assign Y[4'b1111] [35] = 64'h00000000000007A2;
assign u[4'b1111] [35] = 64'h0000000000000BA2;
assign v[4'b1111] [35] = 64'h0000000000000FA2;
assign X[4'b1111] [36] = 64'h00000000000003E3;
assign Y[4'b1111] [36] = 64'h00000000000007A3;
assign u[4'b1111] [36] = 64'h0000000000000BA3;
assign v[4'b1111] [36] = 64'h0000000000000FA3;
assign X[4'b1111] [37] = 64'h00000000000003E4;
assign Y[4'b1111] [37] = 64'h00000000000007A4;
assign u[4'b1111] [37] = 64'h0000000000000BA4;
assign v[4'b1111] [37] = 64'h0000000000000FA4;
assign X[4'b1111] [38] = 64'h00000000000003E5;
assign Y[4'b1111] [38] = 64'h00000000000007A5;
assign u[4'b1111] [38] = 64'h0000000000000BA5;
assign v[4'b1111] [38] = 64'h0000000000000FA5;
assign X[4'b1111] [39] = 64'h00000000000003E6;
assign Y[4'b1111] [39] = 64'h00000000000007A6;
assign u[4'b1111] [39] = 64'h0000000000000BA6;
assign v[4'b1111] [39] = 64'h0000000000000FA6;
assign X[4'b1111] [40] = 64'h00000000000003E7;
assign Y[4'b1111] [40] = 64'h00000000000007A7;
assign u[4'b1111] [40] = 64'h0000000000000BA7;
assign v[4'b1111] [40] = 64'h0000000000000FA7;
assign X[4'b1111] [41] = 64'h00000000000003E8;
assign Y[4'b1111] [41] = 64'h00000000000007A8;
assign u[4'b1111] [41] = 64'h0000000000000BA8;
assign v[4'b1111] [41] = 64'h0000000000000FA8;
assign X[4'b1111] [42] = 64'h00000000000003E9;
assign Y[4'b1111] [42] = 64'h00000000000007A9;
assign u[4'b1111] [42] = 64'h0000000000000BA9;
assign v[4'b1111] [42] = 64'h0000000000000FA9;
assign X[4'b1111] [43] = 64'h00000000000003EA;
assign Y[4'b1111] [43] = 64'h00000000000007AA;
assign u[4'b1111] [43] = 64'h0000000000000BAA;
assign v[4'b1111] [43] = 64'h0000000000000FAA;
assign X[4'b1111] [44] = 64'h00000000000003EB;
assign Y[4'b1111] [44] = 64'h00000000000007AB;
assign u[4'b1111] [44] = 64'h0000000000000BAB;
assign v[4'b1111] [44] = 64'h0000000000000FAB;
assign X[4'b1111] [45] = 64'h00000000000003EC;
assign Y[4'b1111] [45] = 64'h00000000000007AC;
assign u[4'b1111] [45] = 64'h0000000000000BAC;
assign v[4'b1111] [45] = 64'h0000000000000FAC;
assign X[4'b1111] [46] = 64'h00000000000003ED;
assign Y[4'b1111] [46] = 64'h00000000000007AD;
assign u[4'b1111] [46] = 64'h0000000000000BAD;
assign v[4'b1111] [46] = 64'h0000000000000FAD;
assign X[4'b1111] [47] = 64'h00000000000003EE;
assign Y[4'b1111] [47] = 64'h00000000000007AE;
assign u[4'b1111] [47] = 64'h0000000000000BAE;
assign v[4'b1111] [47] = 64'h0000000000000FAE;
assign X[4'b1111] [48] = 64'h00000000000003EF;
assign Y[4'b1111] [48] = 64'h00000000000007AF;
assign u[4'b1111] [48] = 64'h0000000000000BAF;
assign v[4'b1111] [48] = 64'h0000000000000FAF;
assign X[4'b1111] [49] = 64'h00000000000003F0;
assign Y[4'b1111] [49] = 64'h00000000000007B0;
assign u[4'b1111] [49] = 64'h0000000000000BB0;
assign v[4'b1111] [49] = 64'h0000000000000FB0;
assign X[4'b1111] [50] = 64'h00000000000003F1;
assign Y[4'b1111] [50] = 64'h00000000000007B1;
assign u[4'b1111] [50] = 64'h0000000000000BB1;
assign v[4'b1111] [50] = 64'h0000000000000FB1;
assign X[4'b1111] [51] = 64'h00000000000003F2;
assign Y[4'b1111] [51] = 64'h00000000000007B2;
assign u[4'b1111] [51] = 64'h0000000000000BB2;
assign v[4'b1111] [51] = 64'h0000000000000FB2;
assign X[4'b1111] [52] = 64'h00000000000003F3;
assign Y[4'b1111] [52] = 64'h00000000000007B3;
assign u[4'b1111] [52] = 64'h0000000000000BB3;
assign v[4'b1111] [52] = 64'h0000000000000FB3;
assign X[4'b1111] [53] = 64'h00000000000003F4;
assign Y[4'b1111] [53] = 64'h00000000000007B4;
assign u[4'b1111] [53] = 64'h0000000000000BB4;
assign v[4'b1111] [53] = 64'h0000000000000FB4;
assign X[4'b1111] [54] = 64'h00000000000003F5;
assign Y[4'b1111] [54] = 64'h00000000000007B5;
assign u[4'b1111] [54] = 64'h0000000000000BB5;
assign v[4'b1111] [54] = 64'h0000000000000FB5;
assign X[4'b1111] [55] = 64'h00000000000003F6;
assign Y[4'b1111] [55] = 64'h00000000000007B6;
assign u[4'b1111] [55] = 64'h0000000000000BB6;
assign v[4'b1111] [55] = 64'h0000000000000FB6;
assign X[4'b1111] [56] = 64'h00000000000003F7;
assign Y[4'b1111] [56] = 64'h00000000000007B7;
assign u[4'b1111] [56] = 64'h0000000000000BB7;
assign v[4'b1111] [56] = 64'h0000000000000FB7;
assign X[4'b1111] [57] = 64'h00000000000003F8;
assign Y[4'b1111] [57] = 64'h00000000000007B8;
assign u[4'b1111] [57] = 64'h0000000000000BB8;
assign v[4'b1111] [57] = 64'h0000000000000FB8;
assign X[4'b1111] [58] = 64'h00000000000003F9;
assign Y[4'b1111] [58] = 64'h00000000000007B9;
assign u[4'b1111] [58] = 64'h0000000000000BB9;
assign v[4'b1111] [58] = 64'h0000000000000FB9;
assign X[4'b1111] [59] = 64'h00000000000003FA;
assign Y[4'b1111] [59] = 64'h00000000000007BA;
assign u[4'b1111] [59] = 64'h0000000000000BBA;
assign v[4'b1111] [59] = 64'h0000000000000FBA;
assign X[4'b1111] [60] = 64'h00000000000003FB;
assign Y[4'b1111] [60] = 64'h00000000000007BB;
assign u[4'b1111] [60] = 64'h0000000000000BBB;
assign v[4'b1111] [60] = 64'h0000000000000FBB;
assign X[4'b1111] [61] = 64'h00000000000003FC;
assign Y[4'b1111] [61] = 64'h00000000000007BC;
assign u[4'b1111] [61] = 64'h0000000000000BBC;
assign v[4'b1111] [61] = 64'h0000000000000FBC;
assign X[4'b1111] [62] = 64'h00000000000003FD;
assign Y[4'b1111] [62] = 64'h00000000000007BD;
assign u[4'b1111] [62] = 64'h0000000000000BBD;
assign v[4'b1111] [62] = 64'h0000000000000FBD;
assign X[4'b1111] [63] = 64'h00000000000003FE;
assign Y[4'b1111] [63] = 64'h00000000000007BE;
assign u[4'b1111] [63] = 64'h0000000000000BBE;
assign v[4'b1111] [63] = 64'h0000000000000FBE;
assign X[4'b1111] [64] = 64'h00000000000003FF;
assign Y[4'b1111] [64] = 64'h00000000000007BF;
assign u[4'b1111] [64] = 64'h0000000000000BBF;
assign v[4'b1111] [64] = 64'h0000000000000FBF;
