// -----------------------------------------------------------------------------
//
// -----------------------------------------------------------------------------
// Description:
// ------------
//
// Redundant Binary Representation (RBR) adder
//
// Digit |  Value interpreted
// ------|-------------------
// 00    | -1
// 01    |  0
// 10    |  0
// 11    |  1
//
//
// -----------------------------------------------------------------------------
// File name:
// ----------
//
// rbr_add.v
//
// -----------------------------------------------------------------------------
// Interface:
// ----------
//
//  Data inputs:
//    - a         : Summand a (RBR, 2*W bits).
//    - b         : Summand b (RBR, 2*W bits).
//
//  Data outputs:
//    - c         : Result c=a+b (RBR, 2*W bits).
//
//  Parameters:
//    - W         : Word width (natural, default: 64).
//
// -----------------------------------------------------------------------------
// History:
// --------
//
//    - 2016-04-08 - ilesser - Original version.
//
// -----------------------------------------------------------------------------

// *****************************************************************************
// Interface
// *****************************************************************************
module rbr_add #(
    // ----------------------------------
    // Parameters
    // ----------------------------------
    parameter W      = 64
  ) (
    // ----------------------------------
    // Data inputs
    // ----------------------------------
    input   reg   [2*W-1:0]   a,
    input   reg   [2*W-1:0]   b,
    // ----------------------------------
    // Data outputs
    // ----------------------------------
    output  reg   [2*W-1:0]   s,
  );
// *****************************************************************************

// *****************************************************************************
// Architecture
// *****************************************************************************

   // -----------------------------------------------------
   // Internal signals
   // -----------------------------------------------------
   wire [2*W-1:0] c;
   reg  [W-1:0]   sa;
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Combinational logic
   // -----------------------------------------------------
   initial
      c[1]  = 1'b1;
      c[0]  = 1'b0;

   genvar i;
   generate
      for (i=0; i < W-1; i=i+1) begin
         always @(*) begin

            {c[2*(i+1)+1], sa[i]}      = a[2*i+1]  + a[2*i] + b[2*i+1];

            {c[2*(i+1)  ], s[2*i+1]}   = sa[i]     + b[2*i] + c[2*i+1];

            s[2*i] = c[2*i];

         end
      end
   endgenerate
   // -----------------------------------------------------
   // Digit-by-digit diagram
   // -----------------------------------------------------
   //                   a           b
   //                    i           i
   //                   | |         | |
   //                   | |         | |
   //                 +-----+       | |
   //                 |     |       | |
   //           +-----| FA  |-------+ |
   //           |     |     |         |
   //           |     +-----+         |
   //           |        |            |
   //           |     sa | +----------+
   //           |       i| |
   //           |      +-----+
   //           |      |     |
   //   c    ---+   +--| FA  |-----------c
   //    i+1 -------+  |     |       +--- i
   //                  +-----+       |
   //                     |          |
   //                     |+---------+
   //                     ||
   //                     ||
   //                     s
   //                      i
   //
   // -----------------------------------------------------

// *****************************************************************************

// *****************************************************************************
// Assertions and debugging
// *****************************************************************************
`ifdef RTL_DEBUG

   XXXXX TO FILL IN HERE XXXXX

`endif
// *****************************************************************************

endmodule

