assign X[4'b0000] [01] = +0.0000000000000000;
assign Y[4'b0000] [01] = +0.0000000000000000;
assign u[4'b0000] [01] = +0.0000000000000000;
assign v[4'b0000] [01] = +0.0000000000000000;
assign X[4'b0000] [02] = +0.0000000000000000;
assign Y[4'b0000] [02] = +0.0000000000000000;
assign u[4'b0000] [02] = +0.0000000000000000;
assign v[4'b0000] [02] = +0.0000000000000000;
assign X[4'b0000] [03] = +0.0000000000000000;
assign Y[4'b0000] [03] = +0.0000000000000000;
assign u[4'b0000] [03] = +0.0000000000000000;
assign v[4'b0000] [03] = +0.0000000000000000;
assign X[4'b0000] [04] = +0.0000000000000000;
assign Y[4'b0000] [04] = +0.0000000000000000;
assign u[4'b0000] [04] = +0.0000000000000000;
assign v[4'b0000] [04] = +0.0000000000000000;
assign X[4'b0000] [05] = +0.0000000000000000;
assign Y[4'b0000] [05] = +0.0000000000000000;
assign u[4'b0000] [05] = +0.0000000000000000;
assign v[4'b0000] [05] = +0.0000000000000000;
assign X[4'b0000] [06] = +0.0000000000000000;
assign Y[4'b0000] [06] = +0.0000000000000000;
assign u[4'b0000] [06] = +0.0000000000000000;
assign v[4'b0000] [06] = +0.0000000000000000;
assign X[4'b0000] [07] = +0.0000000000000000;
assign Y[4'b0000] [07] = +0.0000000000000000;
assign u[4'b0000] [07] = +0.0000000000000000;
assign v[4'b0000] [07] = +0.0000000000000000;
assign X[4'b0000] [08] = +0.0000000000000000;
assign Y[4'b0000] [08] = +0.0000000000000000;
assign u[4'b0000] [08] = +0.0000000000000000;
assign v[4'b0000] [08] = +0.0000000000000000;
assign X[4'b0000] [09] = +0.0000000000000000;
assign Y[4'b0000] [09] = +0.0000000000000000;
assign u[4'b0000] [09] = +0.0000000000000000;
assign v[4'b0000] [09] = +0.0000000000000000;
assign X[4'b0000] [10] = +0.0000000000000000;
assign Y[4'b0000] [10] = +0.0000000000000000;
assign u[4'b0000] [10] = +0.0000000000000000;
assign v[4'b0000] [10] = +0.0000000000000000;
assign X[4'b0000] [11] = +0.0000000000000000;
assign Y[4'b0000] [11] = +0.0000000000000000;
assign u[4'b0000] [11] = +0.0000000000000000;
assign v[4'b0000] [11] = +0.0000000000000000;
assign X[4'b0000] [12] = +0.0000000000000000;
assign Y[4'b0000] [12] = +0.0000000000000000;
assign u[4'b0000] [12] = +0.0000000000000000;
assign v[4'b0000] [12] = +0.0000000000000000;
assign X[4'b0000] [13] = +0.0000000000000000;
assign Y[4'b0000] [13] = +0.0000000000000000;
assign u[4'b0000] [13] = +0.0000000000000000;
assign v[4'b0000] [13] = +0.0000000000000000;
assign X[4'b0000] [14] = +0.0000000000000000;
assign Y[4'b0000] [14] = +0.0000000000000000;
assign u[4'b0000] [14] = +0.0000000000000000;
assign v[4'b0000] [14] = +0.0000000000000000;
assign X[4'b0000] [15] = +0.0000000000000000;
assign Y[4'b0000] [15] = +0.0000000000000000;
assign u[4'b0000] [15] = +0.0000000000000000;
assign v[4'b0000] [15] = +0.0000000000000000;
assign X[4'b0000] [16] = +0.0000000000000000;
assign Y[4'b0000] [16] = +0.0000000000000000;
assign u[4'b0000] [16] = +0.0000000000000000;
assign v[4'b0000] [16] = +0.0000000000000000;
assign X[4'b0000] [17] = +0.0000000000000000;
assign Y[4'b0000] [17] = +0.0000000000000000;
assign u[4'b0000] [17] = +0.0000000000000000;
assign v[4'b0000] [17] = +0.0000000000000000;
assign X[4'b0000] [18] = +0.0000000000000000;
assign Y[4'b0000] [18] = +0.0000000000000000;
assign u[4'b0000] [18] = +0.0000000000000000;
assign v[4'b0000] [18] = +0.0000000000000000;
assign X[4'b0000] [19] = +0.0000000000000000;
assign Y[4'b0000] [19] = +0.0000000000000000;
assign u[4'b0000] [19] = +0.0000000000000000;
assign v[4'b0000] [19] = +0.0000000000000000;
assign X[4'b0000] [20] = +0.0000000000000000;
assign Y[4'b0000] [20] = +0.0000000000000000;
assign u[4'b0000] [20] = +0.0000000000000000;
assign v[4'b0000] [20] = +0.0000000000000000;
assign X[4'b0000] [21] = +0.0000000000000000;
assign Y[4'b0000] [21] = +0.0000000000000000;
assign u[4'b0000] [21] = +0.0000000000000000;
assign v[4'b0000] [21] = +0.0000000000000000;
assign X[4'b0001] [01] = +0.1115717756571049;
assign Y[4'b0001] [01] = +0.4636476090008061;
assign u[4'b0001] [01] = +0.4462871026284197;
assign v[4'b0001] [01] = +1.8545904360032244;
assign X[4'b0001] [02] = +0.0303123109082174;
assign Y[4'b0001] [02] = +0.2449786631268641;
assign u[4'b0001] [02] = +0.2424984872657394;
assign v[4'b0001] [02] = +1.9598293050149131;
assign X[4'b0001] [03] = +0.0077520932679826;
assign Y[4'b0001] [03] = +0.1243549945467614;
assign u[4'b0001] [03] = +0.1240334922877210;
assign v[4'b0001] [03] = +1.9896799127481830;
assign X[4'b0001] [04] = +0.0019493202078287;
assign Y[4'b0001] [04] = +0.0624188099959574;
assign u[4'b0001] [04] = +0.0623782466505195;
assign v[4'b0001] [04] = +1.9974019198706352;
assign X[4'b0001] [05] = +0.0004880429865277;
assign Y[4'b0001] [05] = +0.0312398334302683;
assign u[4'b0001] [05] = +0.0312347511377731;
assign v[4'b0001] [05] = +1.9993493395371698;
assign X[4'b0001] [06] = +0.0001220554137636;
assign Y[4'b0001] [06] = +0.0156237286204768;
assign u[4'b0001] [06] = +0.0156230929617406;
assign v[4'b0001] [06] = +1.9998372634210344;
assign X[4'b0001] [07] = +0.0000305166468403;
assign Y[4'b0001] [07] = +0.0078123410601011;
assign u[4'b0001] [07] = +0.0078122615911219;
assign v[4'b0001] [07] = +1.9999593113858845;
assign X[4'b0001] [08] = +0.0000076293363242;
assign Y[4'b0001] [08] = +0.0039062301319670;
assign u[4'b0001] [08] = +0.0039062201979808;
assign v[4'b0001] [08] = +1.9999898275670895;
assign X[4'b0001] [09] = +0.0000019073449948;
assign Y[4'b0001] [09] = +0.0019531225164788;
assign u[4'b0001] [09] = +0.0019531212747156;
assign v[4'b0001] [09] = +1.9999974568743104;
assign X[4'b0001] [10] = +0.0000004768369308;
assign Y[4'b0001] [10] = +0.0009765621895593;
assign u[4'b0001] [10] = +0.0009765620343389;
assign v[4'b0001] [10] = +1.9999993642174863;
assign X[4'b0001] [11] = +0.0000001192092753;
assign Y[4'b0001] [11] = +0.0004882812111949;
assign u[4'b0001] [11] = +0.0004882811917923;
assign v[4'b0001] [11] = +1.9999998410543034;
assign X[4'b0001] [12] = +0.0000000298023215;
assign Y[4'b0001] [12] = +0.0002441406201494;
assign u[4'b0001] [12] = +0.0002441406177240;
assign v[4'b0001] [12] = +1.9999999602635716;
assign X[4'b0001] [13] = +0.0000000074505806;
assign Y[4'b0001] [13] = +0.0001220703118937;
assign u[4'b0001] [13] = +0.0001220703120453;
assign v[4'b0001] [13] = +1.9999999900658927;
assign X[4'b0001] [14] = +0.0000000018626451;
assign Y[4'b0001] [14] = +0.0000610351561742;
assign u[4'b0001] [14] = +0.0000610351561932;
assign v[4'b0001] [14] = +1.9999999975164731;
assign X[4'b0001] [15] = +0.0000000004656613;
assign Y[4'b0001] [15] = +0.0000305175781155;
assign u[4'b0001] [15] = +0.0000305175781179;
assign v[4'b0001] [15] = +1.9999999993791182;
assign X[4'b0001] [16] = +0.0000000001164153;
assign Y[4'b0001] [16] = +0.0000152587890613;
assign u[4'b0001] [16] = +0.0000152587890616;
assign v[4'b0001] [16] = +1.9999999998447795;
assign X[4'b0001] [17] = +0.0000000000291038;
assign Y[4'b0001] [17] = +0.0000076293945311;
assign u[4'b0001] [17] = +0.0000076293945311;
assign v[4'b0001] [17] = +1.9999999999611948;
assign X[4'b0001] [18] = +0.0000000000072760;
assign Y[4'b0001] [18] = +0.0000038146972656;
assign u[4'b0001] [18] = +0.0000038146972656;
assign v[4'b0001] [18] = +1.9999999999902986;
assign X[4'b0001] [19] = +0.0000000000018190;
assign Y[4'b0001] [19] = +0.0000019073486328;
assign u[4'b0001] [19] = +0.0000019073486328;
assign v[4'b0001] [19] = +1.9999999999975746;
assign X[4'b0001] [20] = +0.0000000000004547;
assign Y[4'b0001] [20] = +0.0000009536743164;
assign u[4'b0001] [20] = +0.0000009536743164;
assign v[4'b0001] [20] = +1.9999999999993936;
assign X[4'b0001] [21] = +0.0000000000001137;
assign Y[4'b0001] [21] = +0.0000004768371582;
assign u[4'b0001] [21] = +0.0000004768371582;
assign v[4'b0001] [21] = +1.9999999999998483;
assign X[4'b0010] [01] = +0.0000000000000000;
assign Y[4'b0010] [01] = +0.0000000000000000;
assign u[4'b0010] [01] = +0.0000000000000000;
assign v[4'b0010] [01] = +0.0000000000000000;
assign X[4'b0010] [02] = +0.0000000000000000;
assign Y[4'b0010] [02] = +0.0000000000000000;
assign u[4'b0010] [02] = +0.0000000000000000;
assign v[4'b0010] [02] = +0.0000000000000000;
assign X[4'b0010] [03] = +0.0000000000000000;
assign Y[4'b0010] [03] = +0.0000000000000000;
assign u[4'b0010] [03] = +0.0000000000000000;
assign v[4'b0010] [03] = +0.0000000000000000;
assign X[4'b0010] [04] = +0.0000000000000000;
assign Y[4'b0010] [04] = +0.0000000000000000;
assign u[4'b0010] [04] = +0.0000000000000000;
assign v[4'b0010] [04] = +0.0000000000000000;
assign X[4'b0010] [05] = +0.0000000000000000;
assign Y[4'b0010] [05] = +0.0000000000000000;
assign u[4'b0010] [05] = +0.0000000000000000;
assign v[4'b0010] [05] = +0.0000000000000000;
assign X[4'b0010] [06] = +0.0000000000000000;
assign Y[4'b0010] [06] = +0.0000000000000000;
assign u[4'b0010] [06] = +0.0000000000000000;
assign v[4'b0010] [06] = +0.0000000000000000;
assign X[4'b0010] [07] = +0.0000000000000000;
assign Y[4'b0010] [07] = +0.0000000000000000;
assign u[4'b0010] [07] = +0.0000000000000000;
assign v[4'b0010] [07] = +0.0000000000000000;
assign X[4'b0010] [08] = +0.0000000000000000;
assign Y[4'b0010] [08] = +0.0000000000000000;
assign u[4'b0010] [08] = +0.0000000000000000;
assign v[4'b0010] [08] = +0.0000000000000000;
assign X[4'b0010] [09] = +0.0000000000000000;
assign Y[4'b0010] [09] = +0.0000000000000000;
assign u[4'b0010] [09] = +0.0000000000000000;
assign v[4'b0010] [09] = +0.0000000000000000;
assign X[4'b0010] [10] = +0.0000000000000000;
assign Y[4'b0010] [10] = +0.0000000000000000;
assign u[4'b0010] [10] = +0.0000000000000000;
assign v[4'b0010] [10] = +0.0000000000000000;
assign X[4'b0010] [11] = +0.0000000000000000;
assign Y[4'b0010] [11] = +0.0000000000000000;
assign u[4'b0010] [11] = +0.0000000000000000;
assign v[4'b0010] [11] = +0.0000000000000000;
assign X[4'b0010] [12] = +0.0000000000000000;
assign Y[4'b0010] [12] = +0.0000000000000000;
assign u[4'b0010] [12] = +0.0000000000000000;
assign v[4'b0010] [12] = +0.0000000000000000;
assign X[4'b0010] [13] = +0.0000000000000000;
assign Y[4'b0010] [13] = +0.0000000000000000;
assign u[4'b0010] [13] = +0.0000000000000000;
assign v[4'b0010] [13] = +0.0000000000000000;
assign X[4'b0010] [14] = +0.0000000000000000;
assign Y[4'b0010] [14] = +0.0000000000000000;
assign u[4'b0010] [14] = +0.0000000000000000;
assign v[4'b0010] [14] = +0.0000000000000000;
assign X[4'b0010] [15] = +0.0000000000000000;
assign Y[4'b0010] [15] = +0.0000000000000000;
assign u[4'b0010] [15] = +0.0000000000000000;
assign v[4'b0010] [15] = +0.0000000000000000;
assign X[4'b0010] [16] = +0.0000000000000000;
assign Y[4'b0010] [16] = +0.0000000000000000;
assign u[4'b0010] [16] = +0.0000000000000000;
assign v[4'b0010] [16] = +0.0000000000000000;
assign X[4'b0010] [17] = +0.0000000000000000;
assign Y[4'b0010] [17] = +0.0000000000000000;
assign u[4'b0010] [17] = +0.0000000000000000;
assign v[4'b0010] [17] = +0.0000000000000000;
assign X[4'b0010] [18] = +0.0000000000000000;
assign Y[4'b0010] [18] = +0.0000000000000000;
assign u[4'b0010] [18] = +0.0000000000000000;
assign v[4'b0010] [18] = +0.0000000000000000;
assign X[4'b0010] [19] = +0.0000000000000000;
assign Y[4'b0010] [19] = +0.0000000000000000;
assign u[4'b0010] [19] = +0.0000000000000000;
assign v[4'b0010] [19] = +0.0000000000000000;
assign X[4'b0010] [20] = +0.0000000000000000;
assign Y[4'b0010] [20] = +0.0000000000000000;
assign u[4'b0010] [20] = +0.0000000000000000;
assign v[4'b0010] [20] = +0.0000000000000000;
assign X[4'b0010] [21] = +0.0000000000000000;
assign Y[4'b0010] [21] = +0.0000000000000000;
assign u[4'b0010] [21] = +0.0000000000000000;
assign v[4'b0010] [21] = +0.0000000000000000;
assign X[4'b0011] [01] = +0.1115717756571049;
assign Y[4'b0011] [01] = -0.4636476090008061;
assign u[4'b0011] [01] = +0.4462871026284197;
assign v[4'b0011] [01] = -1.8545904360032244;
assign X[4'b0011] [02] = +0.0303123109082174;
assign Y[4'b0011] [02] = -0.2449786631268641;
assign u[4'b0011] [02] = +0.2424984872657394;
assign v[4'b0011] [02] = -1.9598293050149131;
assign X[4'b0011] [03] = +0.0077520932679826;
assign Y[4'b0011] [03] = -0.1243549945467614;
assign u[4'b0011] [03] = +0.1240334922877210;
assign v[4'b0011] [03] = -1.9896799127481830;
assign X[4'b0011] [04] = +0.0019493202078287;
assign Y[4'b0011] [04] = -0.0624188099959574;
assign u[4'b0011] [04] = +0.0623782466505195;
assign v[4'b0011] [04] = -1.9974019198706352;
assign X[4'b0011] [05] = +0.0004880429865277;
assign Y[4'b0011] [05] = -0.0312398334302683;
assign u[4'b0011] [05] = +0.0312347511377731;
assign v[4'b0011] [05] = -1.9993493395371698;
assign X[4'b0011] [06] = +0.0001220554137636;
assign Y[4'b0011] [06] = -0.0156237286204768;
assign u[4'b0011] [06] = +0.0156230929617406;
assign v[4'b0011] [06] = -1.9998372634210344;
assign X[4'b0011] [07] = +0.0000305166468403;
assign Y[4'b0011] [07] = -0.0078123410601011;
assign u[4'b0011] [07] = +0.0078122615911219;
assign v[4'b0011] [07] = -1.9999593113858845;
assign X[4'b0011] [08] = +0.0000076293363242;
assign Y[4'b0011] [08] = -0.0039062301319670;
assign u[4'b0011] [08] = +0.0039062201979808;
assign v[4'b0011] [08] = -1.9999898275670895;
assign X[4'b0011] [09] = +0.0000019073449948;
assign Y[4'b0011] [09] = -0.0019531225164788;
assign u[4'b0011] [09] = +0.0019531212747156;
assign v[4'b0011] [09] = -1.9999974568743104;
assign X[4'b0011] [10] = +0.0000004768369308;
assign Y[4'b0011] [10] = -0.0009765621895593;
assign u[4'b0011] [10] = +0.0009765620343389;
assign v[4'b0011] [10] = -1.9999993642174863;
assign X[4'b0011] [11] = +0.0000001192092753;
assign Y[4'b0011] [11] = -0.0004882812111949;
assign u[4'b0011] [11] = +0.0004882811917923;
assign v[4'b0011] [11] = -1.9999998410543034;
assign X[4'b0011] [12] = +0.0000000298023215;
assign Y[4'b0011] [12] = -0.0002441406201494;
assign u[4'b0011] [12] = +0.0002441406177240;
assign v[4'b0011] [12] = -1.9999999602635716;
assign X[4'b0011] [13] = +0.0000000074505806;
assign Y[4'b0011] [13] = -0.0001220703118937;
assign u[4'b0011] [13] = +0.0001220703120453;
assign v[4'b0011] [13] = -1.9999999900658927;
assign X[4'b0011] [14] = +0.0000000018626451;
assign Y[4'b0011] [14] = -0.0000610351561742;
assign u[4'b0011] [14] = +0.0000610351561932;
assign v[4'b0011] [14] = -1.9999999975164731;
assign X[4'b0011] [15] = +0.0000000004656613;
assign Y[4'b0011] [15] = -0.0000305175781155;
assign u[4'b0011] [15] = +0.0000305175781179;
assign v[4'b0011] [15] = -1.9999999993791182;
assign X[4'b0011] [16] = +0.0000000001164153;
assign Y[4'b0011] [16] = -0.0000152587890613;
assign u[4'b0011] [16] = +0.0000152587890616;
assign v[4'b0011] [16] = -1.9999999998447795;
assign X[4'b0011] [17] = +0.0000000000291038;
assign Y[4'b0011] [17] = -0.0000076293945311;
assign u[4'b0011] [17] = +0.0000076293945311;
assign v[4'b0011] [17] = -1.9999999999611948;
assign X[4'b0011] [18] = +0.0000000000072760;
assign Y[4'b0011] [18] = -0.0000038146972656;
assign u[4'b0011] [18] = +0.0000038146972656;
assign v[4'b0011] [18] = -1.9999999999902986;
assign X[4'b0011] [19] = +0.0000000000018190;
assign Y[4'b0011] [19] = -0.0000019073486328;
assign u[4'b0011] [19] = +0.0000019073486328;
assign v[4'b0011] [19] = -1.9999999999975746;
assign X[4'b0011] [20] = +0.0000000000004547;
assign Y[4'b0011] [20] = -0.0000009536743164;
assign u[4'b0011] [20] = +0.0000009536743164;
assign v[4'b0011] [20] = -1.9999999999993936;
assign X[4'b0011] [21] = +0.0000000000001137;
assign Y[4'b0011] [21] = -0.0000004768371582;
assign u[4'b0011] [21] = +0.0000004768371582;
assign v[4'b0011] [21] = -1.9999999999998483;
assign X[4'b0100] [01] = +0.4054651081081644;
assign Y[4'b0100] [01] = +0.0000000000000000;
assign u[4'b0100] [01] = +1.6218604324326575;
assign v[4'b0100] [01] = +0.0000000000000000;
assign X[4'b0100] [02] = +0.2231435513142098;
assign Y[4'b0100] [02] = +0.0000000000000000;
assign u[4'b0100] [02] = +1.7851484105136781;
assign v[4'b0100] [02] = +0.0000000000000000;
assign X[4'b0100] [03] = +0.1177830356563835;
assign Y[4'b0100] [03] = +0.0000000000000000;
assign u[4'b0100] [03] = +1.8845285705021353;
assign v[4'b0100] [03] = +0.0000000000000000;
assign X[4'b0100] [04] = +0.0606246218164348;
assign Y[4'b0100] [04] = +0.0000000000000000;
assign u[4'b0100] [04] = +1.9399878981259149;
assign v[4'b0100] [04] = +0.0000000000000000;
assign X[4'b0100] [05] = +0.0307716586667537;
assign Y[4'b0100] [05] = +0.0000000000000000;
assign u[4'b0100] [05] = +1.9693861546722360;
assign v[4'b0100] [05] = +0.0000000000000000;
assign X[4'b0100] [06] = +0.0155041865359653;
assign Y[4'b0100] [06] = +0.0000000000000000;
assign u[4'b0100] [06] = +1.9845358766035526;
assign v[4'b0100] [06] = +0.0000000000000000;
assign X[4'b0100] [07] = +0.0077821404420549;
assign Y[4'b0100] [07] = +0.0000000000000000;
assign u[4'b0100] [07] = +1.9922279531660669;
assign v[4'b0100] [07] = +0.0000000000000000;
assign X[4'b0100] [08] = +0.0038986404156573;
assign Y[4'b0100] [08] = +0.0000000000000000;
assign u[4'b0100] [08] = +1.9961038928165493;
assign v[4'b0100] [08] = +0.0000000000000000;
assign X[4'b0100] [09] = +0.0019512201312617;
assign Y[4'b0100] [09] = +0.0000000000000000;
assign u[4'b0100] [09] = +1.9980494144120313;
assign v[4'b0100] [09] = +0.0000000000000000;
assign X[4'b0100] [10] = +0.0009760859730555;
assign Y[4'b0100] [10] = +0.0000000000000000;
assign u[4'b0100] [10] = +1.9990240728175799;
assign v[4'b0100] [10] = +0.0000000000000000;
assign X[4'b0100] [11] = +0.0004881620795014;
assign Y[4'b0100] [11] = +0.0000000000000000;
assign u[4'b0100] [11] = +1.9995118776375345;
assign v[4'b0100] [11] = +0.0000000000000000;
assign X[4'b0100] [12] = +0.0002441108275274;
assign Y[4'b0100] [12] = +0.0000000000000000;
assign u[4'b0100] [12] = +1.9997558991041553;
assign v[4'b0100] [12] = +0.0000000000000000;
assign X[4'b0100] [13] = +0.0001220628625257;
assign Y[4'b0100] [13] = +0.0000000000000000;
assign u[4'b0100] [13] = +1.9998779396206980;
assign v[4'b0100] [13] = +0.0000000000000000;
assign X[4'b0100] [14] = +0.0000610332936806;
assign Y[4'b0100] [14] = +0.0000000000000000;
assign u[4'b0100] [14] = +1.9999389673271633;
assign v[4'b0100] [14] = +0.0000000000000000;
assign X[4'b0100] [15] = +0.0000305171124732;
assign Y[4'b0100] [15] = +0.0000000000000000;
assign u[4'b0100] [15] = +1.9999694830427426;
assign v[4'b0100] [15] = +0.0000000000000000;
assign X[4'b0100] [16] = +0.0000152586726484;
assign Y[4'b0100] [16] = +0.0000000000000000;
assign u[4'b0100] [16] = +1.9999847413661562;
assign v[4'b0100] [16] = +0.0000000000000000;
assign X[4'b0100] [17] = +0.0000076293654276;
assign Y[4'b0100] [17] = +0.0000000000000000;
assign u[4'b0100] [17] = +1.9999923706442737;
assign v[4'b0100] [17] = +0.0000000000000000;
assign X[4'b0100] [18] = +0.0000038146899897;
assign Y[4'b0100] [18] = +0.0000000000000000;
assign u[4'b0100] [18] = +1.9999961853124357;
assign v[4'b0100] [18] = +0.0000000000000000;
assign X[4'b0100] [19] = +0.0000019073468138;
assign Y[4'b0100] [19] = +0.0000000000000000;
assign u[4'b0100] [19] = +1.9999980926537926;
assign v[4'b0100] [19] = +0.0000000000000000;
assign X[4'b0100] [20] = +0.0000009536738617;
assign Y[4'b0100] [20] = +0.0000000000000000;
assign u[4'b0100] [20] = +1.9999990463262900;
assign v[4'b0100] [20] = +0.0000000000000000;
assign X[4'b0100] [21] = +0.0000004768370445;
assign Y[4'b0100] [21] = +0.0000000000000000;
assign u[4'b0100] [21] = +1.9999995231629935;
assign v[4'b0100] [21] = +0.0000000000000000;
assign X[4'b0101] [01] = +0.4581453659370776;
assign Y[4'b0101] [01] = +0.3217505543966422;
assign u[4'b0101] [01] = +1.8325814637483104;
assign v[4'b0101] [01] = +1.2870022175865687;
assign X[4'b0101] [02] = +0.2427539078908503;
assign Y[4'b0101] [02] = +0.1973955598498807;
assign u[4'b0101] [02] = +1.9420312631268026;
assign v[4'b0101] [02] = +1.5791644787990460;
assign X[4'b0101] [03] = +0.1239180819522907;
assign Y[4'b0101] [03] = +0.1106572211738956;
assign u[4'b0101] [03] = +1.9826893112366513;
assign v[4'b0101] [03] = +1.7705155387823304;
assign X[4'b0101] [04] = +0.0623517392504787;
assign Y[4'b0101] [04] = +0.0587558227157227;
assign u[4'b0101] [04] = +1.9952556560153185;
assign v[4'b0101] [04] = +1.8801863269031263;
assign X[4'b0101] [05] = +0.0312305848118681;
assign Y[4'b0101] [05] = +0.0302937599187751;
assign u[4'b0101] [05] = +1.9987574279595595;
assign v[4'b0101] [05] = +1.9388006348016065;
assign X[4'b0101] [06] = +0.0156225157283291;
assign Y[4'b0101] [06] = +0.0153834017805952;
assign u[4'b0101] [06] = +1.9996820132261188;
assign v[4'b0101] [06] = +1.9690754279161793;
assign X[4'b0101] [07] = +0.0078121858105703;
assign Y[4'b0101] [07] = +0.0077517827122069;
assign u[4'b0101] [07] = +1.9999195675060046;
assign v[4'b0101] [07] = +1.9844563743249595;
assign X[4'b0101] [08] = +0.0039062104956732;
assign Y[4'b0101] [08] = +0.0038910309466445;
assign u[4'b0101] [08] = +1.9999797737846823;
assign v[4'b0101] [08] = +1.9922078446819715;
assign X[4'b0101] [09] = +0.0019531200474755;
assign Y[4'b0101] [09] = +0.0019493152697654;
assign u[4'b0101] [09] = +1.9999949286148679;
assign v[4'b0101] [09] = +1.9960988362398133;
assign X[4'b0101] [10] = +0.0009765618800270;
assign Y[4'b0101] [10] = +0.0009756094465646;
assign u[4'b0101] [10] = +1.9999987302952080;
assign v[4'b0101] [10] = +1.9980481465643023;
assign X[4'b0101] [11] = +0.0004882811724466;
assign Y[4'b0101] [11] = +0.0004880429090311;
assign u[4'b0101] [11] = +1.9999996823413151;
assign v[4'b0101] [11] = +1.9990237553913479;
assign X[4'b0101] [12] = +0.0002441406153023;
assign Y[4'b0101] [12] = +0.0002440810300565;
assign u[4'b0101] [12] = +1.9999999205562393;
assign v[4'b0101] [12] = +1.9995117982228541;
assign X[4'b0101] [13] = +0.0001220703112875;
assign Y[4'b0101] [13] = +0.0001220554125515;
assign u[4'b0101] [13] = +1.9999999801340587;
assign v[4'b0101] [13] = +1.9997558792432146;
assign X[4'b0101] [14] = +0.0000610351560984;
assign Y[4'b0101] [14] = +0.0000610314311113;
assign u[4'b0101] [14] = +1.9999999950332306;
assign v[4'b0101] [14] = +1.9998779346545537;
assign X[4'b0101] [15] = +0.0000305175781061;
assign Y[4'b0101] [15] = +0.0000305166468214;
assign u[4'b0101] [15] = +1.9999999987582722;
assign v[4'b0101] [15] = +1.9999389660855134;
assign X[4'b0101] [16] = +0.0000152587890601;
assign Y[4'b0101] [16] = +0.0000152585562342;
assign u[4'b0101] [16] = +1.9999999996895637;
assign v[4'b0101] [16] = +1.9999694827323158;
assign X[4'b0101] [17] = +0.0000076293945310;
assign Y[4'b0101] [17] = +0.0000076293363239;
assign u[4'b0101] [17] = +1.9999999999223903;
assign v[4'b0101] [17] = +1.9999847412885476;
assign X[4'b0101] [18] = +0.0000038146972656;
assign Y[4'b0101] [18] = +0.0000038146827137;
assign u[4'b0101] [18] = +1.9999999999951494;
assign v[4'b0101] [18] = +1.9999923706248712;
assign X[4'b0101] [19] = +0.0000019073486328;
assign Y[4'b0101] [19] = +0.0000019073449948;
assign u[4'b0101] [19] = +1.9999999999987874;
assign v[4'b0101] [19] = +1.9999961853075849;
assign X[4'b0101] [20] = +0.0000009536743164;
assign Y[4'b0101] [20] = +0.0000009536734069;
assign u[4'b0101] [20] = +1.9999999999996969;
assign v[4'b0101] [20] = +1.9999980926525798;
assign X[4'b0101] [21] = +0.0000004768371582;
assign Y[4'b0101] [21] = +0.0000004768369308;
assign u[4'b0101] [21] = +1.9999999999999243;
assign v[4'b0101] [21] = +1.9999990463259867;
assign X[4'b0110] [01] = +0.4054651081081644;
assign Y[4'b0110] [01] = +0.0000000000000000;
assign u[4'b0110] [01] = +1.6218604324326575;
assign v[4'b0110] [01] = +0.0000000000000000;
assign X[4'b0110] [02] = +0.2231435513142098;
assign Y[4'b0110] [02] = +0.0000000000000000;
assign u[4'b0110] [02] = +1.7851484105136781;
assign v[4'b0110] [02] = +0.0000000000000000;
assign X[4'b0110] [03] = +0.1177830356563835;
assign Y[4'b0110] [03] = +0.0000000000000000;
assign u[4'b0110] [03] = +1.8845285705021353;
assign v[4'b0110] [03] = +0.0000000000000000;
assign X[4'b0110] [04] = +0.0606246218164348;
assign Y[4'b0110] [04] = +0.0000000000000000;
assign u[4'b0110] [04] = +1.9399878981259149;
assign v[4'b0110] [04] = +0.0000000000000000;
assign X[4'b0110] [05] = +0.0307716586667537;
assign Y[4'b0110] [05] = +0.0000000000000000;
assign u[4'b0110] [05] = +1.9693861546722360;
assign v[4'b0110] [05] = +0.0000000000000000;
assign X[4'b0110] [06] = +0.0155041865359653;
assign Y[4'b0110] [06] = +0.0000000000000000;
assign u[4'b0110] [06] = +1.9845358766035526;
assign v[4'b0110] [06] = +0.0000000000000000;
assign X[4'b0110] [07] = +0.0077821404420549;
assign Y[4'b0110] [07] = +0.0000000000000000;
assign u[4'b0110] [07] = +1.9922279531660669;
assign v[4'b0110] [07] = +0.0000000000000000;
assign X[4'b0110] [08] = +0.0038986404156573;
assign Y[4'b0110] [08] = +0.0000000000000000;
assign u[4'b0110] [08] = +1.9961038928165493;
assign v[4'b0110] [08] = +0.0000000000000000;
assign X[4'b0110] [09] = +0.0019512201312617;
assign Y[4'b0110] [09] = +0.0000000000000000;
assign u[4'b0110] [09] = +1.9980494144120313;
assign v[4'b0110] [09] = +0.0000000000000000;
assign X[4'b0110] [10] = +0.0009760859730555;
assign Y[4'b0110] [10] = +0.0000000000000000;
assign u[4'b0110] [10] = +1.9990240728175799;
assign v[4'b0110] [10] = +0.0000000000000000;
assign X[4'b0110] [11] = +0.0004881620795014;
assign Y[4'b0110] [11] = +0.0000000000000000;
assign u[4'b0110] [11] = +1.9995118776375345;
assign v[4'b0110] [11] = +0.0000000000000000;
assign X[4'b0110] [12] = +0.0002441108275274;
assign Y[4'b0110] [12] = +0.0000000000000000;
assign u[4'b0110] [12] = +1.9997558991041553;
assign v[4'b0110] [12] = +0.0000000000000000;
assign X[4'b0110] [13] = +0.0001220628625257;
assign Y[4'b0110] [13] = +0.0000000000000000;
assign u[4'b0110] [13] = +1.9998779396206980;
assign v[4'b0110] [13] = +0.0000000000000000;
assign X[4'b0110] [14] = +0.0000610332936806;
assign Y[4'b0110] [14] = +0.0000000000000000;
assign u[4'b0110] [14] = +1.9999389673271633;
assign v[4'b0110] [14] = +0.0000000000000000;
assign X[4'b0110] [15] = +0.0000305171124732;
assign Y[4'b0110] [15] = +0.0000000000000000;
assign u[4'b0110] [15] = +1.9999694830427426;
assign v[4'b0110] [15] = +0.0000000000000000;
assign X[4'b0110] [16] = +0.0000152586726484;
assign Y[4'b0110] [16] = +0.0000000000000000;
assign u[4'b0110] [16] = +1.9999847413661562;
assign v[4'b0110] [16] = +0.0000000000000000;
assign X[4'b0110] [17] = +0.0000076293654276;
assign Y[4'b0110] [17] = +0.0000000000000000;
assign u[4'b0110] [17] = +1.9999923706442737;
assign v[4'b0110] [17] = +0.0000000000000000;
assign X[4'b0110] [18] = +0.0000038146899897;
assign Y[4'b0110] [18] = +0.0000000000000000;
assign u[4'b0110] [18] = +1.9999961853124357;
assign v[4'b0110] [18] = +0.0000000000000000;
assign X[4'b0110] [19] = +0.0000019073468138;
assign Y[4'b0110] [19] = +0.0000000000000000;
assign u[4'b0110] [19] = +1.9999980926537926;
assign v[4'b0110] [19] = +0.0000000000000000;
assign X[4'b0110] [20] = +0.0000009536738617;
assign Y[4'b0110] [20] = +0.0000000000000000;
assign u[4'b0110] [20] = +1.9999990463262900;
assign v[4'b0110] [20] = +0.0000000000000000;
assign X[4'b0110] [21] = +0.0000004768370445;
assign Y[4'b0110] [21] = +0.0000000000000000;
assign u[4'b0110] [21] = +1.9999995231629935;
assign v[4'b0110] [21] = +0.0000000000000000;
assign X[4'b0111] [01] = +0.4581453659370776;
assign Y[4'b0111] [01] = -0.3217505543966422;
assign u[4'b0111] [01] = +1.8325814637483104;
assign v[4'b0111] [01] = -1.2870022175865687;
assign X[4'b0111] [02] = +0.2427539078908503;
assign Y[4'b0111] [02] = -0.1973955598498807;
assign u[4'b0111] [02] = +1.9420312631268026;
assign v[4'b0111] [02] = -1.5791644787990460;
assign X[4'b0111] [03] = +0.1239180819522907;
assign Y[4'b0111] [03] = -0.1106572211738956;
assign u[4'b0111] [03] = +1.9826893112366513;
assign v[4'b0111] [03] = -1.7705155387823304;
assign X[4'b0111] [04] = +0.0623517392504787;
assign Y[4'b0111] [04] = -0.0587558227157227;
assign u[4'b0111] [04] = +1.9952556560153185;
assign v[4'b0111] [04] = -1.8801863269031263;
assign X[4'b0111] [05] = +0.0312305848118681;
assign Y[4'b0111] [05] = -0.0302937599187751;
assign u[4'b0111] [05] = +1.9987574279595595;
assign v[4'b0111] [05] = -1.9388006348016065;
assign X[4'b0111] [06] = +0.0156225157283291;
assign Y[4'b0111] [06] = -0.0153834017805952;
assign u[4'b0111] [06] = +1.9996820132261188;
assign v[4'b0111] [06] = -1.9690754279161793;
assign X[4'b0111] [07] = +0.0078121858105703;
assign Y[4'b0111] [07] = -0.0077517827122069;
assign u[4'b0111] [07] = +1.9999195675060046;
assign v[4'b0111] [07] = -1.9844563743249595;
assign X[4'b0111] [08] = +0.0039062104956732;
assign Y[4'b0111] [08] = -0.0038910309466445;
assign u[4'b0111] [08] = +1.9999797737846823;
assign v[4'b0111] [08] = -1.9922078446819715;
assign X[4'b0111] [09] = +0.0019531200474755;
assign Y[4'b0111] [09] = -0.0019493152697654;
assign u[4'b0111] [09] = +1.9999949286148679;
assign v[4'b0111] [09] = -1.9960988362398133;
assign X[4'b0111] [10] = +0.0009765618800270;
assign Y[4'b0111] [10] = -0.0009756094465646;
assign u[4'b0111] [10] = +1.9999987302952080;
assign v[4'b0111] [10] = -1.9980481465643023;
assign X[4'b0111] [11] = +0.0004882811724466;
assign Y[4'b0111] [11] = -0.0004880429090311;
assign u[4'b0111] [11] = +1.9999996823413151;
assign v[4'b0111] [11] = -1.9990237553913479;
assign X[4'b0111] [12] = +0.0002441406153023;
assign Y[4'b0111] [12] = -0.0002440810300565;
assign u[4'b0111] [12] = +1.9999999205562393;
assign v[4'b0111] [12] = -1.9995117982228541;
assign X[4'b0111] [13] = +0.0001220703112875;
assign Y[4'b0111] [13] = -0.0001220554125515;
assign u[4'b0111] [13] = +1.9999999801340587;
assign v[4'b0111] [13] = -1.9997558792432146;
assign X[4'b0111] [14] = +0.0000610351560984;
assign Y[4'b0111] [14] = -0.0000610314311113;
assign u[4'b0111] [14] = +1.9999999950332306;
assign v[4'b0111] [14] = -1.9998779346545537;
assign X[4'b0111] [15] = +0.0000305175781061;
assign Y[4'b0111] [15] = -0.0000305166468214;
assign u[4'b0111] [15] = +1.9999999987582722;
assign v[4'b0111] [15] = -1.9999389660855134;
assign X[4'b0111] [16] = +0.0000152587890601;
assign Y[4'b0111] [16] = -0.0000152585562342;
assign u[4'b0111] [16] = +1.9999999996895637;
assign v[4'b0111] [16] = -1.9999694827323158;
assign X[4'b0111] [17] = +0.0000076293945310;
assign Y[4'b0111] [17] = -0.0000076293363239;
assign u[4'b0111] [17] = +1.9999999999223903;
assign v[4'b0111] [17] = -1.9999847412885476;
assign X[4'b0111] [18] = +0.0000038146972656;
assign Y[4'b0111] [18] = -0.0000038146827137;
assign u[4'b0111] [18] = +1.9999999999951494;
assign v[4'b0111] [18] = -1.9999923706248712;
assign X[4'b0111] [19] = +0.0000019073486328;
assign Y[4'b0111] [19] = -0.0000019073449948;
assign u[4'b0111] [19] = +1.9999999999987874;
assign v[4'b0111] [19] = -1.9999961853075849;
assign X[4'b0111] [20] = +0.0000009536743164;
assign Y[4'b0111] [20] = -0.0000009536734069;
assign u[4'b0111] [20] = +1.9999999999996969;
assign v[4'b0111] [20] = -1.9999980926525798;
assign X[4'b0111] [21] = +0.0000004768371582;
assign Y[4'b0111] [21] = -0.0000004768369308;
assign u[4'b0111] [21] = +1.9999999999999243;
assign v[4'b0111] [21] = -1.9999990463259867;
assign X[4'b1000] [01] = +0.0000000000000000;
assign Y[4'b1000] [01] = +0.0000000000000000;
assign u[4'b1000] [01] = +0.0000000000000000;
assign v[4'b1000] [01] = +0.0000000000000000;
assign X[4'b1000] [02] = +0.0000000000000000;
assign Y[4'b1000] [02] = +0.0000000000000000;
assign u[4'b1000] [02] = +0.0000000000000000;
assign v[4'b1000] [02] = +0.0000000000000000;
assign X[4'b1000] [03] = +0.0000000000000000;
assign Y[4'b1000] [03] = +0.0000000000000000;
assign u[4'b1000] [03] = +0.0000000000000000;
assign v[4'b1000] [03] = +0.0000000000000000;
assign X[4'b1000] [04] = +0.0000000000000000;
assign Y[4'b1000] [04] = +0.0000000000000000;
assign u[4'b1000] [04] = +0.0000000000000000;
assign v[4'b1000] [04] = +0.0000000000000000;
assign X[4'b1000] [05] = +0.0000000000000000;
assign Y[4'b1000] [05] = +0.0000000000000000;
assign u[4'b1000] [05] = +0.0000000000000000;
assign v[4'b1000] [05] = +0.0000000000000000;
assign X[4'b1000] [06] = +0.0000000000000000;
assign Y[4'b1000] [06] = +0.0000000000000000;
assign u[4'b1000] [06] = +0.0000000000000000;
assign v[4'b1000] [06] = +0.0000000000000000;
assign X[4'b1000] [07] = +0.0000000000000000;
assign Y[4'b1000] [07] = +0.0000000000000000;
assign u[4'b1000] [07] = +0.0000000000000000;
assign v[4'b1000] [07] = +0.0000000000000000;
assign X[4'b1000] [08] = +0.0000000000000000;
assign Y[4'b1000] [08] = +0.0000000000000000;
assign u[4'b1000] [08] = +0.0000000000000000;
assign v[4'b1000] [08] = +0.0000000000000000;
assign X[4'b1000] [09] = +0.0000000000000000;
assign Y[4'b1000] [09] = +0.0000000000000000;
assign u[4'b1000] [09] = +0.0000000000000000;
assign v[4'b1000] [09] = +0.0000000000000000;
assign X[4'b1000] [10] = +0.0000000000000000;
assign Y[4'b1000] [10] = +0.0000000000000000;
assign u[4'b1000] [10] = +0.0000000000000000;
assign v[4'b1000] [10] = +0.0000000000000000;
assign X[4'b1000] [11] = +0.0000000000000000;
assign Y[4'b1000] [11] = +0.0000000000000000;
assign u[4'b1000] [11] = +0.0000000000000000;
assign v[4'b1000] [11] = +0.0000000000000000;
assign X[4'b1000] [12] = +0.0000000000000000;
assign Y[4'b1000] [12] = +0.0000000000000000;
assign u[4'b1000] [12] = +0.0000000000000000;
assign v[4'b1000] [12] = +0.0000000000000000;
assign X[4'b1000] [13] = +0.0000000000000000;
assign Y[4'b1000] [13] = +0.0000000000000000;
assign u[4'b1000] [13] = +0.0000000000000000;
assign v[4'b1000] [13] = +0.0000000000000000;
assign X[4'b1000] [14] = +0.0000000000000000;
assign Y[4'b1000] [14] = +0.0000000000000000;
assign u[4'b1000] [14] = +0.0000000000000000;
assign v[4'b1000] [14] = +0.0000000000000000;
assign X[4'b1000] [15] = +0.0000000000000000;
assign Y[4'b1000] [15] = +0.0000000000000000;
assign u[4'b1000] [15] = +0.0000000000000000;
assign v[4'b1000] [15] = +0.0000000000000000;
assign X[4'b1000] [16] = +0.0000000000000000;
assign Y[4'b1000] [16] = +0.0000000000000000;
assign u[4'b1000] [16] = +0.0000000000000000;
assign v[4'b1000] [16] = +0.0000000000000000;
assign X[4'b1000] [17] = +0.0000000000000000;
assign Y[4'b1000] [17] = +0.0000000000000000;
assign u[4'b1000] [17] = +0.0000000000000000;
assign v[4'b1000] [17] = +0.0000000000000000;
assign X[4'b1000] [18] = +0.0000000000000000;
assign Y[4'b1000] [18] = +0.0000000000000000;
assign u[4'b1000] [18] = +0.0000000000000000;
assign v[4'b1000] [18] = +0.0000000000000000;
assign X[4'b1000] [19] = +0.0000000000000000;
assign Y[4'b1000] [19] = +0.0000000000000000;
assign u[4'b1000] [19] = +0.0000000000000000;
assign v[4'b1000] [19] = +0.0000000000000000;
assign X[4'b1000] [20] = +0.0000000000000000;
assign Y[4'b1000] [20] = +0.0000000000000000;
assign u[4'b1000] [20] = +0.0000000000000000;
assign v[4'b1000] [20] = +0.0000000000000000;
assign X[4'b1000] [21] = +0.0000000000000000;
assign Y[4'b1000] [21] = +0.0000000000000000;
assign u[4'b1000] [21] = +0.0000000000000000;
assign v[4'b1000] [21] = +0.0000000000000000;
assign X[4'b1001] [01] = +0.1115717756571049;
assign Y[4'b1001] [01] = +0.4636476090008061;
assign u[4'b1001] [01] = +0.4462871026284197;
assign v[4'b1001] [01] = +1.8545904360032244;
assign X[4'b1001] [02] = +0.0303123109082174;
assign Y[4'b1001] [02] = +0.2449786631268641;
assign u[4'b1001] [02] = +0.2424984872657394;
assign v[4'b1001] [02] = +1.9598293050149131;
assign X[4'b1001] [03] = +0.0077520932679826;
assign Y[4'b1001] [03] = +0.1243549945467614;
assign u[4'b1001] [03] = +0.1240334922877210;
assign v[4'b1001] [03] = +1.9896799127481830;
assign X[4'b1001] [04] = +0.0019493202078287;
assign Y[4'b1001] [04] = +0.0624188099959574;
assign u[4'b1001] [04] = +0.0623782466505195;
assign v[4'b1001] [04] = +1.9974019198706352;
assign X[4'b1001] [05] = +0.0004880429865277;
assign Y[4'b1001] [05] = +0.0312398334302683;
assign u[4'b1001] [05] = +0.0312347511377731;
assign v[4'b1001] [05] = +1.9993493395371698;
assign X[4'b1001] [06] = +0.0001220554137636;
assign Y[4'b1001] [06] = +0.0156237286204768;
assign u[4'b1001] [06] = +0.0156230929617406;
assign v[4'b1001] [06] = +1.9998372634210344;
assign X[4'b1001] [07] = +0.0000305166468403;
assign Y[4'b1001] [07] = +0.0078123410601011;
assign u[4'b1001] [07] = +0.0078122615911219;
assign v[4'b1001] [07] = +1.9999593113858845;
assign X[4'b1001] [08] = +0.0000076293363242;
assign Y[4'b1001] [08] = +0.0039062301319670;
assign u[4'b1001] [08] = +0.0039062201979808;
assign v[4'b1001] [08] = +1.9999898275670895;
assign X[4'b1001] [09] = +0.0000019073449948;
assign Y[4'b1001] [09] = +0.0019531225164788;
assign u[4'b1001] [09] = +0.0019531212747156;
assign v[4'b1001] [09] = +1.9999974568743104;
assign X[4'b1001] [10] = +0.0000004768369308;
assign Y[4'b1001] [10] = +0.0009765621895593;
assign u[4'b1001] [10] = +0.0009765620343389;
assign v[4'b1001] [10] = +1.9999993642174863;
assign X[4'b1001] [11] = +0.0000001192092753;
assign Y[4'b1001] [11] = +0.0004882812111949;
assign u[4'b1001] [11] = +0.0004882811917923;
assign v[4'b1001] [11] = +1.9999998410543034;
assign X[4'b1001] [12] = +0.0000000298023215;
assign Y[4'b1001] [12] = +0.0002441406201494;
assign u[4'b1001] [12] = +0.0002441406177240;
assign v[4'b1001] [12] = +1.9999999602635716;
assign X[4'b1001] [13] = +0.0000000074505806;
assign Y[4'b1001] [13] = +0.0001220703118937;
assign u[4'b1001] [13] = +0.0001220703120453;
assign v[4'b1001] [13] = +1.9999999900658927;
assign X[4'b1001] [14] = +0.0000000018626451;
assign Y[4'b1001] [14] = +0.0000610351561742;
assign u[4'b1001] [14] = +0.0000610351561932;
assign v[4'b1001] [14] = +1.9999999975164731;
assign X[4'b1001] [15] = +0.0000000004656613;
assign Y[4'b1001] [15] = +0.0000305175781155;
assign u[4'b1001] [15] = +0.0000305175781179;
assign v[4'b1001] [15] = +1.9999999993791182;
assign X[4'b1001] [16] = +0.0000000001164153;
assign Y[4'b1001] [16] = +0.0000152587890613;
assign u[4'b1001] [16] = +0.0000152587890616;
assign v[4'b1001] [16] = +1.9999999998447795;
assign X[4'b1001] [17] = +0.0000000000291038;
assign Y[4'b1001] [17] = +0.0000076293945311;
assign u[4'b1001] [17] = +0.0000076293945311;
assign v[4'b1001] [17] = +1.9999999999611948;
assign X[4'b1001] [18] = +0.0000000000072760;
assign Y[4'b1001] [18] = +0.0000038146972656;
assign u[4'b1001] [18] = +0.0000038146972656;
assign v[4'b1001] [18] = +1.9999999999902986;
assign X[4'b1001] [19] = +0.0000000000018190;
assign Y[4'b1001] [19] = +0.0000019073486328;
assign u[4'b1001] [19] = +0.0000019073486328;
assign v[4'b1001] [19] = +1.9999999999975746;
assign X[4'b1001] [20] = +0.0000000000004547;
assign Y[4'b1001] [20] = +0.0000009536743164;
assign u[4'b1001] [20] = +0.0000009536743164;
assign v[4'b1001] [20] = +1.9999999999993936;
assign X[4'b1001] [21] = +0.0000000000001137;
assign Y[4'b1001] [21] = +0.0000004768371582;
assign u[4'b1001] [21] = +0.0000004768371582;
assign v[4'b1001] [21] = +1.9999999999998483;
assign X[4'b1010] [01] = +0.0000000000000000;
assign Y[4'b1010] [01] = +0.0000000000000000;
assign u[4'b1010] [01] = +0.0000000000000000;
assign v[4'b1010] [01] = +0.0000000000000000;
assign X[4'b1010] [02] = +0.0000000000000000;
assign Y[4'b1010] [02] = +0.0000000000000000;
assign u[4'b1010] [02] = +0.0000000000000000;
assign v[4'b1010] [02] = +0.0000000000000000;
assign X[4'b1010] [03] = +0.0000000000000000;
assign Y[4'b1010] [03] = +0.0000000000000000;
assign u[4'b1010] [03] = +0.0000000000000000;
assign v[4'b1010] [03] = +0.0000000000000000;
assign X[4'b1010] [04] = +0.0000000000000000;
assign Y[4'b1010] [04] = +0.0000000000000000;
assign u[4'b1010] [04] = +0.0000000000000000;
assign v[4'b1010] [04] = +0.0000000000000000;
assign X[4'b1010] [05] = +0.0000000000000000;
assign Y[4'b1010] [05] = +0.0000000000000000;
assign u[4'b1010] [05] = +0.0000000000000000;
assign v[4'b1010] [05] = +0.0000000000000000;
assign X[4'b1010] [06] = +0.0000000000000000;
assign Y[4'b1010] [06] = +0.0000000000000000;
assign u[4'b1010] [06] = +0.0000000000000000;
assign v[4'b1010] [06] = +0.0000000000000000;
assign X[4'b1010] [07] = +0.0000000000000000;
assign Y[4'b1010] [07] = +0.0000000000000000;
assign u[4'b1010] [07] = +0.0000000000000000;
assign v[4'b1010] [07] = +0.0000000000000000;
assign X[4'b1010] [08] = +0.0000000000000000;
assign Y[4'b1010] [08] = +0.0000000000000000;
assign u[4'b1010] [08] = +0.0000000000000000;
assign v[4'b1010] [08] = +0.0000000000000000;
assign X[4'b1010] [09] = +0.0000000000000000;
assign Y[4'b1010] [09] = +0.0000000000000000;
assign u[4'b1010] [09] = +0.0000000000000000;
assign v[4'b1010] [09] = +0.0000000000000000;
assign X[4'b1010] [10] = +0.0000000000000000;
assign Y[4'b1010] [10] = +0.0000000000000000;
assign u[4'b1010] [10] = +0.0000000000000000;
assign v[4'b1010] [10] = +0.0000000000000000;
assign X[4'b1010] [11] = +0.0000000000000000;
assign Y[4'b1010] [11] = +0.0000000000000000;
assign u[4'b1010] [11] = +0.0000000000000000;
assign v[4'b1010] [11] = +0.0000000000000000;
assign X[4'b1010] [12] = +0.0000000000000000;
assign Y[4'b1010] [12] = +0.0000000000000000;
assign u[4'b1010] [12] = +0.0000000000000000;
assign v[4'b1010] [12] = +0.0000000000000000;
assign X[4'b1010] [13] = +0.0000000000000000;
assign Y[4'b1010] [13] = +0.0000000000000000;
assign u[4'b1010] [13] = +0.0000000000000000;
assign v[4'b1010] [13] = +0.0000000000000000;
assign X[4'b1010] [14] = +0.0000000000000000;
assign Y[4'b1010] [14] = +0.0000000000000000;
assign u[4'b1010] [14] = +0.0000000000000000;
assign v[4'b1010] [14] = +0.0000000000000000;
assign X[4'b1010] [15] = +0.0000000000000000;
assign Y[4'b1010] [15] = +0.0000000000000000;
assign u[4'b1010] [15] = +0.0000000000000000;
assign v[4'b1010] [15] = +0.0000000000000000;
assign X[4'b1010] [16] = +0.0000000000000000;
assign Y[4'b1010] [16] = +0.0000000000000000;
assign u[4'b1010] [16] = +0.0000000000000000;
assign v[4'b1010] [16] = +0.0000000000000000;
assign X[4'b1010] [17] = +0.0000000000000000;
assign Y[4'b1010] [17] = +0.0000000000000000;
assign u[4'b1010] [17] = +0.0000000000000000;
assign v[4'b1010] [17] = +0.0000000000000000;
assign X[4'b1010] [18] = +0.0000000000000000;
assign Y[4'b1010] [18] = +0.0000000000000000;
assign u[4'b1010] [18] = +0.0000000000000000;
assign v[4'b1010] [18] = +0.0000000000000000;
assign X[4'b1010] [19] = +0.0000000000000000;
assign Y[4'b1010] [19] = +0.0000000000000000;
assign u[4'b1010] [19] = +0.0000000000000000;
assign v[4'b1010] [19] = +0.0000000000000000;
assign X[4'b1010] [20] = +0.0000000000000000;
assign Y[4'b1010] [20] = +0.0000000000000000;
assign u[4'b1010] [20] = +0.0000000000000000;
assign v[4'b1010] [20] = +0.0000000000000000;
assign X[4'b1010] [21] = +0.0000000000000000;
assign Y[4'b1010] [21] = +0.0000000000000000;
assign u[4'b1010] [21] = +0.0000000000000000;
assign v[4'b1010] [21] = +0.0000000000000000;
assign X[4'b1011] [01] = +0.1115717756571049;
assign Y[4'b1011] [01] = -0.4636476090008061;
assign u[4'b1011] [01] = +0.4462871026284197;
assign v[4'b1011] [01] = -1.8545904360032244;
assign X[4'b1011] [02] = +0.0303123109082174;
assign Y[4'b1011] [02] = -0.2449786631268641;
assign u[4'b1011] [02] = +0.2424984872657394;
assign v[4'b1011] [02] = -1.9598293050149131;
assign X[4'b1011] [03] = +0.0077520932679826;
assign Y[4'b1011] [03] = -0.1243549945467614;
assign u[4'b1011] [03] = +0.1240334922877210;
assign v[4'b1011] [03] = -1.9896799127481830;
assign X[4'b1011] [04] = +0.0019493202078287;
assign Y[4'b1011] [04] = -0.0624188099959574;
assign u[4'b1011] [04] = +0.0623782466505195;
assign v[4'b1011] [04] = -1.9974019198706352;
assign X[4'b1011] [05] = +0.0004880429865277;
assign Y[4'b1011] [05] = -0.0312398334302683;
assign u[4'b1011] [05] = +0.0312347511377731;
assign v[4'b1011] [05] = -1.9993493395371698;
assign X[4'b1011] [06] = +0.0001220554137636;
assign Y[4'b1011] [06] = -0.0156237286204768;
assign u[4'b1011] [06] = +0.0156230929617406;
assign v[4'b1011] [06] = -1.9998372634210344;
assign X[4'b1011] [07] = +0.0000305166468403;
assign Y[4'b1011] [07] = -0.0078123410601011;
assign u[4'b1011] [07] = +0.0078122615911219;
assign v[4'b1011] [07] = -1.9999593113858845;
assign X[4'b1011] [08] = +0.0000076293363242;
assign Y[4'b1011] [08] = -0.0039062301319670;
assign u[4'b1011] [08] = +0.0039062201979808;
assign v[4'b1011] [08] = -1.9999898275670895;
assign X[4'b1011] [09] = +0.0000019073449948;
assign Y[4'b1011] [09] = -0.0019531225164788;
assign u[4'b1011] [09] = +0.0019531212747156;
assign v[4'b1011] [09] = -1.9999974568743104;
assign X[4'b1011] [10] = +0.0000004768369308;
assign Y[4'b1011] [10] = -0.0009765621895593;
assign u[4'b1011] [10] = +0.0009765620343389;
assign v[4'b1011] [10] = -1.9999993642174863;
assign X[4'b1011] [11] = +0.0000001192092753;
assign Y[4'b1011] [11] = -0.0004882812111949;
assign u[4'b1011] [11] = +0.0004882811917923;
assign v[4'b1011] [11] = -1.9999998410543034;
assign X[4'b1011] [12] = +0.0000000298023215;
assign Y[4'b1011] [12] = -0.0002441406201494;
assign u[4'b1011] [12] = +0.0002441406177240;
assign v[4'b1011] [12] = -1.9999999602635716;
assign X[4'b1011] [13] = +0.0000000074505806;
assign Y[4'b1011] [13] = -0.0001220703118937;
assign u[4'b1011] [13] = +0.0001220703120453;
assign v[4'b1011] [13] = -1.9999999900658927;
assign X[4'b1011] [14] = +0.0000000018626451;
assign Y[4'b1011] [14] = -0.0000610351561742;
assign u[4'b1011] [14] = +0.0000610351561932;
assign v[4'b1011] [14] = -1.9999999975164731;
assign X[4'b1011] [15] = +0.0000000004656613;
assign Y[4'b1011] [15] = -0.0000305175781155;
assign u[4'b1011] [15] = +0.0000305175781179;
assign v[4'b1011] [15] = -1.9999999993791182;
assign X[4'b1011] [16] = +0.0000000001164153;
assign Y[4'b1011] [16] = -0.0000152587890613;
assign u[4'b1011] [16] = +0.0000152587890616;
assign v[4'b1011] [16] = -1.9999999998447795;
assign X[4'b1011] [17] = +0.0000000000291038;
assign Y[4'b1011] [17] = -0.0000076293945311;
assign u[4'b1011] [17] = +0.0000076293945311;
assign v[4'b1011] [17] = -1.9999999999611948;
assign X[4'b1011] [18] = +0.0000000000072760;
assign Y[4'b1011] [18] = -0.0000038146972656;
assign u[4'b1011] [18] = +0.0000038146972656;
assign v[4'b1011] [18] = -1.9999999999902986;
assign X[4'b1011] [19] = +0.0000000000018190;
assign Y[4'b1011] [19] = -0.0000019073486328;
assign u[4'b1011] [19] = +0.0000019073486328;
assign v[4'b1011] [19] = -1.9999999999975746;
assign X[4'b1011] [20] = +0.0000000000004547;
assign Y[4'b1011] [20] = -0.0000009536743164;
assign u[4'b1011] [20] = +0.0000009536743164;
assign v[4'b1011] [20] = -1.9999999999993936;
assign X[4'b1011] [21] = +0.0000000000001137;
assign Y[4'b1011] [21] = -0.0000004768371582;
assign u[4'b1011] [21] = +0.0000004768371582;
assign v[4'b1011] [21] = -1.9999999999998483;
assign X[4'b1100] [01] = -0.6931471805599453;
assign Y[4'b1100] [01] = +0.0000000000000000;
assign u[4'b1100] [01] = -2.7725887222397811;
assign v[4'b1100] [01] = +0.0000000000000000;
assign X[4'b1100] [02] = -0.2876820724517809;
assign Y[4'b1100] [02] = +0.0000000000000000;
assign u[4'b1100] [02] = -2.3014565796142472;
assign v[4'b1100] [02] = +0.0000000000000000;
assign X[4'b1100] [03] = -0.1335313926245226;
assign Y[4'b1100] [03] = +0.0000000000000000;
assign u[4'b1100] [03] = -2.1365022819923620;
assign v[4'b1100] [03] = +0.0000000000000000;
assign X[4'b1100] [04] = -0.0645385211375712;
assign Y[4'b1100] [04] = +0.0000000000000000;
assign u[4'b1100] [04] = -2.0652326764022777;
assign v[4'b1100] [04] = +0.0000000000000000;
assign X[4'b1100] [05] = -0.0317486983145803;
assign Y[4'b1100] [05] = +0.0000000000000000;
assign u[4'b1100] [05] = -2.0319166921331391;
assign v[4'b1100] [05] = +0.0000000000000000;
assign X[4'b1100] [06] = -0.0157483569681392;
assign Y[4'b1100] [06] = +0.0000000000000000;
assign u[4'b1100] [06] = -2.0157896919218135;
assign v[4'b1100] [06] = +0.0000000000000000;
assign X[4'b1100] [07] = -0.0078431774610259;
assign Y[4'b1100] [07] = +0.0000000000000000;
assign u[4'b1100] [07] = -2.0078534300226285;
assign v[4'b1100] [07] = +0.0000000000000000;
assign X[4'b1100] [08] = -0.0039138993211363;
assign Y[4'b1100] [08] = +0.0000000000000000;
assign u[4'b1100] [08] = -2.0039164524218003;
assign v[4'b1100] [08] = +0.0000000000000000;
assign X[4'b1100] [09] = -0.0019550348358034;
assign Y[4'b1100] [09] = +0.0000000000000000;
assign u[4'b1100] [09] = -2.0019556718626310;
assign v[4'b1100] [09] = +0.0000000000000000;
assign X[4'b1100] [10] = -0.0009770396478266;
assign Y[4'b1100] [10] = +0.0000000000000000;
assign u[4'b1100] [10] = -2.0009771987489029;
assign v[4'b1100] [10] = +0.0000000000000000;
assign X[4'b1100] [11] = -0.0004884004981089;
assign Y[4'b1100] [11] = +0.0000000000000000;
assign u[4'b1100] [11] = -2.0004884402539500;
assign v[4'b1100] [11] = +0.0000000000000000;
assign X[4'b1100] [12] = -0.0002441704321739;
assign Y[4'b1100] [12] = +0.0000000000000000;
assign u[4'b1100] [12] = -2.0002441803687074;
assign v[4'b1100] [12] = +0.0000000000000000;
assign X[4'b1100] [13] = -0.0001220777636870;
assign Y[4'b1100] [13] = +0.0000000000000000;
assign u[4'b1100] [13] = -2.0001220802475173;
assign v[4'b1100] [13] = +0.0000000000000000;
assign X[4'b1100] [14] = -0.0000610370189709;
assign Y[4'b1100] [14] = +0.0000000000000000;
assign u[4'b1100] [14] = -2.0000610376398904;
assign v[4'b1100] [14] = +0.0000000000000000;
assign X[4'b1100] [15] = -0.0000305180437958;
assign Y[4'b1100] [15] = +0.0000000000000000;
assign u[4'b1100] [15] = -2.0000305181990208;
assign v[4'b1100] [15] = +0.0000000000000000;
assign X[4'b1100] [16] = -0.0000152589054790;
assign Y[4'b1100] [16] = +0.0000000000000000;
assign u[4'b1100] [16] = -2.0000152589442846;
assign v[4'b1100] [16] = +0.0000000000000000;
assign X[4'b1100] [17] = -0.0000076294236352;
assign Y[4'b1100] [17] = +0.0000000000000000;
assign u[4'b1100] [17] = -2.0000076294333367;
assign v[4'b1100] [17] = +0.0000000000000000;
assign X[4'b1100] [18] = -0.0000038147045416;
assign Y[4'b1100] [18] = +0.0000000000000000;
assign u[4'b1100] [18] = -2.0000038147069668;
assign v[4'b1100] [18] = +0.0000000000000000;
assign X[4'b1100] [19] = -0.0000019073504518;
assign Y[4'b1100] [19] = +0.0000000000000000;
assign u[4'b1100] [19] = -2.0000019073510580;
assign v[4'b1100] [19] = +0.0000000000000000;
assign X[4'b1100] [20] = -0.0000009536747712;
assign Y[4'b1100] [20] = +0.0000000000000000;
assign u[4'b1100] [20] = -2.0000009536749226;
assign v[4'b1100] [20] = +0.0000000000000000;
assign X[4'b1100] [21] = -0.0000004768372719;
assign Y[4'b1100] [21] = +0.0000000000000000;
assign u[4'b1100] [21] = -2.0000004768373096;
assign v[4'b1100] [21] = +0.0000000000000000;
assign X[4'b1101] [01] = -0.3465735902799726;
assign Y[4'b1101] [01] = +0.7853981633974483;
assign u[4'b1101] [01] = -1.3862943611198904;
assign v[4'b1101] [01] = +3.1415926535897931;
assign X[4'b1101] [02] = -0.2350018146228677;
assign Y[4'b1101] [02] = +0.3217505543966422;
assign u[4'b1101] [02] = -1.8800145169829416;
assign v[4'b1101] [02] = +2.5740044351731375;
assign X[4'b1101] [03] = -0.1234300389657629;
assign Y[4'b1101] [03] = +0.1418970546041639;
assign u[4'b1101] [03] = -1.9748806234522058;
assign v[4'b1101] [03] = +2.2703528736666230;
assign X[4'b1101] [04] = -0.0623212226036383;
assign Y[4'b1101] [04] = +0.0665681637758238;
assign u[4'b1101] [04] = -1.9942791233164259;
assign v[4'b1101] [04] = +2.1301812408263618;
assign X[4'b1101] [05] = -0.0312286774668733;
assign Y[4'b1101] [05] = +0.0322468824352539;
assign u[4'b1101] [05] = -1.9986353578798890;
assign v[4'b1101] [05] = +2.0638004758562509;
assign X[4'b1101] [06] = -0.0156223965190538;
assign Y[4'b1101] [06] = +0.0158716829917901;
assign u[4'b1101] [06] = -1.9996667544388824;
assign v[4'b1101] [06] = +2.0315754229491265;
assign X[4'b1101] [07] = -0.0078121783599899;
assign Y[4'b1101] [07] = +0.0078738530241005;
assign u[4'b1101] [07] = -1.9999176601574109;
assign v[4'b1101] [07] = +2.0157063741697390;
assign X[4'b1101] [08] = -0.0039062100300119;
assign Y[4'b1101] [08] = +0.0039215485247600;
assign u[4'b1101] [08] = -1.9999795353661032;
assign v[4'b1101] [08] = +2.0078328446771208;
assign X[4'b1101] [09] = -0.0019531200183716;
assign Y[4'b1101] [09] = +0.0019569446642965;
assign u[4'b1101] [09] = -1.9999948988125242;
assign v[4'b1101] [09] = +2.0039113362396619;
assign X[4'b1101] [10] = -0.0009765618782081;
assign Y[4'b1101] [10] = +0.0009775167951974;
assign u[4'b1101] [10] = -1.9999987265701442;
assign v[4'b1101] [10] = +2.0019543965642979;
assign X[4'b1101] [11] = -0.0004882811723329;
assign Y[4'b1101] [11] = +0.0004885197461893;
assign u[4'b1101] [11] = -1.9999996818756538;
assign v[4'b1101] [11] = +2.0009768803913479;
assign X[4'b1101] [12] = -0.0002441406152952;
assign Y[4'b1101] [12] = +0.0002442002393461;
assign u[4'b1101] [12] = -1.9999999204980317;
assign v[4'b1101] [12] = +2.0004883607228541;
assign X[4'b1101] [13] = -0.0001220703112871;
assign Y[4'b1101] [13] = +0.0001220852148739;
assign u[4'b1101] [13] = -1.9999999801276920;
assign v[4'b1101] [13] = +2.0002441604932146;
assign X[4'b1101] [14] = -0.0000610351560984;
assign Y[4'b1101] [14] = +0.0000610388816919;
assign u[4'b1101] [14] = -1.9999999950326621;
assign v[4'b1101] [14] = +2.0001220752795539;
assign X[4'b1101] [15] = -0.0000305175781061;
assign Y[4'b1101] [15] = +0.0000305185094665;
assign u[4'b1101] [15] = -1.9999999987582011;
assign v[4'b1101] [15] = +2.0000610363980136;
assign X[4'b1101] [16] = -0.0000152587890601;
assign Y[4'b1101] [16] = +0.0000152590218955;
assign u[4'b1101] [16] = -1.9999999996895548;
assign v[4'b1101] [16] = +2.0000305178885660;
assign X[4'b1101] [17] = -0.0000076293945310;
assign Y[4'b1101] [17] = +0.0000076294527392;
assign u[4'b1101] [17] = -1.9999999999223892;
assign v[4'b1101] [17] = +2.0000152588666729;
assign X[4'b1101] [18] = -0.0000038146972656;
assign Y[4'b1101] [18] = +0.0000038147118176;
assign u[4'b1101] [18] = -1.9999999999951494;
assign v[4'b1101] [18] = +2.0000076294139340;
assign X[4'b1101] [19] = -0.0000019073486328;
assign Y[4'b1101] [19] = +0.0000019073522708;
assign u[4'b1101] [19] = -1.9999999999987874;
assign v[4'b1101] [19] = +2.0000038147021164;
assign X[4'b1101] [20] = -0.0000009536743164;
assign Y[4'b1101] [20] = +0.0000009536752259;
assign u[4'b1101] [20] = -1.9999999999996969;
assign v[4'b1101] [20] = +2.0000019073498456;
assign X[4'b1101] [21] = -0.0000004768371582;
assign Y[4'b1101] [21] = +0.0000004768373856;
assign u[4'b1101] [21] = -1.9999999999999243;
assign v[4'b1101] [21] = +2.0000009536746197;
assign X[4'b1110] [01] = -0.6931471805599453;
assign Y[4'b1110] [01] = +0.0000000000000000;
assign u[4'b1110] [01] = -2.7725887222397811;
assign v[4'b1110] [01] = +0.0000000000000000;
assign X[4'b1110] [02] = -0.2876820724517809;
assign Y[4'b1110] [02] = +0.0000000000000000;
assign u[4'b1110] [02] = -2.3014565796142472;
assign v[4'b1110] [02] = +0.0000000000000000;
assign X[4'b1110] [03] = -0.1335313926245226;
assign Y[4'b1110] [03] = +0.0000000000000000;
assign u[4'b1110] [03] = -2.1365022819923620;
assign v[4'b1110] [03] = +0.0000000000000000;
assign X[4'b1110] [04] = -0.0645385211375712;
assign Y[4'b1110] [04] = +0.0000000000000000;
assign u[4'b1110] [04] = -2.0652326764022777;
assign v[4'b1110] [04] = +0.0000000000000000;
assign X[4'b1110] [05] = -0.0317486983145803;
assign Y[4'b1110] [05] = +0.0000000000000000;
assign u[4'b1110] [05] = -2.0319166921331391;
assign v[4'b1110] [05] = +0.0000000000000000;
assign X[4'b1110] [06] = -0.0157483569681392;
assign Y[4'b1110] [06] = +0.0000000000000000;
assign u[4'b1110] [06] = -2.0157896919218135;
assign v[4'b1110] [06] = +0.0000000000000000;
assign X[4'b1110] [07] = -0.0078431774610259;
assign Y[4'b1110] [07] = +0.0000000000000000;
assign u[4'b1110] [07] = -2.0078534300226285;
assign v[4'b1110] [07] = +0.0000000000000000;
assign X[4'b1110] [08] = -0.0039138993211363;
assign Y[4'b1110] [08] = +0.0000000000000000;
assign u[4'b1110] [08] = -2.0039164524218003;
assign v[4'b1110] [08] = +0.0000000000000000;
assign X[4'b1110] [09] = -0.0019550348358034;
assign Y[4'b1110] [09] = +0.0000000000000000;
assign u[4'b1110] [09] = -2.0019556718626310;
assign v[4'b1110] [09] = +0.0000000000000000;
assign X[4'b1110] [10] = -0.0009770396478266;
assign Y[4'b1110] [10] = +0.0000000000000000;
assign u[4'b1110] [10] = -2.0009771987489029;
assign v[4'b1110] [10] = +0.0000000000000000;
assign X[4'b1110] [11] = -0.0004884004981089;
assign Y[4'b1110] [11] = +0.0000000000000000;
assign u[4'b1110] [11] = -2.0004884402539500;
assign v[4'b1110] [11] = +0.0000000000000000;
assign X[4'b1110] [12] = -0.0002441704321739;
assign Y[4'b1110] [12] = +0.0000000000000000;
assign u[4'b1110] [12] = -2.0002441803687074;
assign v[4'b1110] [12] = +0.0000000000000000;
assign X[4'b1110] [13] = -0.0001220777636870;
assign Y[4'b1110] [13] = +0.0000000000000000;
assign u[4'b1110] [13] = -2.0001220802475173;
assign v[4'b1110] [13] = +0.0000000000000000;
assign X[4'b1110] [14] = -0.0000610370189709;
assign Y[4'b1110] [14] = +0.0000000000000000;
assign u[4'b1110] [14] = -2.0000610376398904;
assign v[4'b1110] [14] = +0.0000000000000000;
assign X[4'b1110] [15] = -0.0000305180437958;
assign Y[4'b1110] [15] = +0.0000000000000000;
assign u[4'b1110] [15] = -2.0000305181990208;
assign v[4'b1110] [15] = +0.0000000000000000;
assign X[4'b1110] [16] = -0.0000152589054790;
assign Y[4'b1110] [16] = +0.0000000000000000;
assign u[4'b1110] [16] = -2.0000152589442846;
assign v[4'b1110] [16] = +0.0000000000000000;
assign X[4'b1110] [17] = -0.0000076294236352;
assign Y[4'b1110] [17] = +0.0000000000000000;
assign u[4'b1110] [17] = -2.0000076294333367;
assign v[4'b1110] [17] = +0.0000000000000000;
assign X[4'b1110] [18] = -0.0000038147045416;
assign Y[4'b1110] [18] = +0.0000000000000000;
assign u[4'b1110] [18] = -2.0000038147069668;
assign v[4'b1110] [18] = +0.0000000000000000;
assign X[4'b1110] [19] = -0.0000019073504518;
assign Y[4'b1110] [19] = +0.0000000000000000;
assign u[4'b1110] [19] = -2.0000019073510580;
assign v[4'b1110] [19] = +0.0000000000000000;
assign X[4'b1110] [20] = -0.0000009536747712;
assign Y[4'b1110] [20] = +0.0000000000000000;
assign u[4'b1110] [20] = -2.0000009536749226;
assign v[4'b1110] [20] = +0.0000000000000000;
assign X[4'b1110] [21] = -0.0000004768372719;
assign Y[4'b1110] [21] = +0.0000000000000000;
assign u[4'b1110] [21] = -2.0000004768373096;
assign v[4'b1110] [21] = +0.0000000000000000;
assign X[4'b1111] [01] = -0.3465735902799726;
assign Y[4'b1111] [01] = -0.7853981633974483;
assign u[4'b1111] [01] = -1.3862943611198904;
assign v[4'b1111] [01] = -3.1415926535897931;
assign X[4'b1111] [02] = -0.2350018146228677;
assign Y[4'b1111] [02] = -0.3217505543966422;
assign u[4'b1111] [02] = -1.8800145169829416;
assign v[4'b1111] [02] = -2.5740044351731375;
assign X[4'b1111] [03] = -0.1234300389657629;
assign Y[4'b1111] [03] = -0.1418970546041639;
assign u[4'b1111] [03] = -1.9748806234522058;
assign v[4'b1111] [03] = -2.2703528736666230;
assign X[4'b1111] [04] = -0.0623212226036383;
assign Y[4'b1111] [04] = -0.0665681637758238;
assign u[4'b1111] [04] = -1.9942791233164259;
assign v[4'b1111] [04] = -2.1301812408263618;
assign X[4'b1111] [05] = -0.0312286774668733;
assign Y[4'b1111] [05] = -0.0322468824352539;
assign u[4'b1111] [05] = -1.9986353578798890;
assign v[4'b1111] [05] = -2.0638004758562509;
assign X[4'b1111] [06] = -0.0156223965190538;
assign Y[4'b1111] [06] = -0.0158716829917901;
assign u[4'b1111] [06] = -1.9996667544388824;
assign v[4'b1111] [06] = -2.0315754229491265;
assign X[4'b1111] [07] = -0.0078121783599899;
assign Y[4'b1111] [07] = -0.0078738530241005;
assign u[4'b1111] [07] = -1.9999176601574109;
assign v[4'b1111] [07] = -2.0157063741697390;
assign X[4'b1111] [08] = -0.0039062100300119;
assign Y[4'b1111] [08] = -0.0039215485247600;
assign u[4'b1111] [08] = -1.9999795353661032;
assign v[4'b1111] [08] = -2.0078328446771208;
assign X[4'b1111] [09] = -0.0019531200183716;
assign Y[4'b1111] [09] = -0.0019569446642965;
assign u[4'b1111] [09] = -1.9999948988125242;
assign v[4'b1111] [09] = -2.0039113362396619;
assign X[4'b1111] [10] = -0.0009765618782081;
assign Y[4'b1111] [10] = -0.0009775167951974;
assign u[4'b1111] [10] = -1.9999987265701442;
assign v[4'b1111] [10] = -2.0019543965642979;
assign X[4'b1111] [11] = -0.0004882811723329;
assign Y[4'b1111] [11] = -0.0004885197461893;
assign u[4'b1111] [11] = -1.9999996818756538;
assign v[4'b1111] [11] = -2.0009768803913479;
assign X[4'b1111] [12] = -0.0002441406152952;
assign Y[4'b1111] [12] = -0.0002442002393461;
assign u[4'b1111] [12] = -1.9999999204980317;
assign v[4'b1111] [12] = -2.0004883607228541;
assign X[4'b1111] [13] = -0.0001220703112871;
assign Y[4'b1111] [13] = -0.0001220852148739;
assign u[4'b1111] [13] = -1.9999999801276920;
assign v[4'b1111] [13] = -2.0002441604932146;
assign X[4'b1111] [14] = -0.0000610351560984;
assign Y[4'b1111] [14] = -0.0000610388816919;
assign u[4'b1111] [14] = -1.9999999950326621;
assign v[4'b1111] [14] = -2.0001220752795539;
assign X[4'b1111] [15] = -0.0000305175781061;
assign Y[4'b1111] [15] = -0.0000305185094665;
assign u[4'b1111] [15] = -1.9999999987582011;
assign v[4'b1111] [15] = -2.0000610363980136;
assign X[4'b1111] [16] = -0.0000152587890601;
assign Y[4'b1111] [16] = -0.0000152590218955;
assign u[4'b1111] [16] = -1.9999999996895548;
assign v[4'b1111] [16] = -2.0000305178885660;
assign X[4'b1111] [17] = -0.0000076293945310;
assign Y[4'b1111] [17] = -0.0000076294527392;
assign u[4'b1111] [17] = -1.9999999999223892;
assign v[4'b1111] [17] = -2.0000152588666729;
assign X[4'b1111] [18] = -0.0000038146972656;
assign Y[4'b1111] [18] = -0.0000038147118176;
assign u[4'b1111] [18] = -1.9999999999951494;
assign v[4'b1111] [18] = -2.0000076294139340;
assign X[4'b1111] [19] = -0.0000019073486328;
assign Y[4'b1111] [19] = -0.0000019073522708;
assign u[4'b1111] [19] = -1.9999999999987874;
assign v[4'b1111] [19] = -2.0000038147021164;
assign X[4'b1111] [20] = -0.0000009536743164;
assign Y[4'b1111] [20] = -0.0000009536752259;
assign u[4'b1111] [20] = -1.9999999999996969;
assign v[4'b1111] [20] = -2.0000019073498456;
assign X[4'b1111] [21] = -0.0000004768371582;
assign Y[4'b1111] [21] = -0.0000004768373856;
assign u[4'b1111] [21] = -1.9999999999999243;
assign v[4'b1111] [21] = -2.0000009536746197;
