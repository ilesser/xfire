// -----------------------------------------------------------------------------
//
// -----------------------------------------------------------------------------
// Description:
// ------------
//
// XXXXX FILL IN HERE XXXXX
//
// -----------------------------------------------------------------------------
// File name:
// ----------
//
// output_precision_selection.v
//
// -----------------------------------------------------------------------------
// Interface:
// ----------
//
//  Clock, reset & enable inputs:
//    - clk      : Posedge active clock input (logic, 1 bit).
//    - arst     : High active asynchronous reset (logic, 1 bit).
//    - enable   : Synchronous enable (logic, 1 bit).
//    - srst     : High active synchronous reset (logic, 1 bit).
//
//  Data inputs:
//    - XXXXX    : XXXXXXXXXX (XXXXX, XXXX bits).
//
//  Data outputs:
//    - XXXXX    : XXXXXXXXXX (XXXXX, XXXX bits).
//
//  Parameters:
//    - XXXXX    : XXXXXXXXXX (XXXXX, default: XXXXX).
//
// -----------------------------------------------------------------------------
// History:
// --------
//
//    - 2016-04-20 - ilesser - Original version.
//
// -----------------------------------------------------------------------------

`include "XXXXXXXX.vh"

// *****************************************************************************
// Interface
// *****************************************************************************
module output_precision_selection #(
    // ----------------------------------
    // Parameters
    // ----------------------------------
    parameter W      = 64
  ) (
    // ----------------------------------
    // Data inputs
    // ----------------------------------
    input wire  [W-1:0]       X_in,
    input wire  [W-1:0]       X_in,
    // ----------------------------------
    // Data outputs
    // ----------------------------------
    output reg  [W-1:0]       X_out,
    output reg  [W-1:0]       X_out
  );
// *****************************************************************************

// *****************************************************************************
// Architecture
// *****************************************************************************

   // -----------------------------------------------------
   // Internal signals
   // -----------------------------------------------------
   // -----------------------------------------------------

   always @(*) begin
      case (format)
         FORMAT_REAL_32:
                        begin
                           X_out = {{W/2{X_in[W/2-1]}},X_in};
                           Y_out = {W{1'b0}};
                        end
         FORMAT_REAL_64:
                        begin
                           X_out = X_in;
                           Y_out = {W{1'b0}};
                        end
         FORMAT_CMPLX_32:
                        begin
                           X_out = {{W/2{X_in[W/2-1]}},X_in};
                           Y_out = {{W/2{Y_in[W/2-1]}},Y_in};
                        end
         FORMAT_CMPLX_64:
                        begin
                           X_out = X_in;
                           Y_out = Y_in;
                        end
         default:
                        begin
                           X_out = {W{1'b0}};
                           Y_out = {W{1'b0}};
                        end
      endcase
   end

// *****************************************************************************

// *****************************************************************************
// Assertions and debugging
// *****************************************************************************
`ifdef RTL_DEBUG

   //XXXXX TO FILL IN HERE XXXXX

`endif
// *****************************************************************************

endmodule

