// -----------------------------------------------------------------------------
//  Copyright (c) 2016 Microelectronics Lab. FIUBA.
//  All Rights Reserved.
//
//  The information contained in this file is confidential and proprietary.
//  Any reproduction, use or disclosure, in whole or in part, of this
//  program, including any attempt to obtain a human-readable version of this
//  program, without the express, prior written consent of Microelectronics Lab.
//  FIUBA is strictly prohibited.
//
// -----------------------------------------------------------------------------
// Description:
// ------------
//
// XXXXX FILL IN HERE XXXXX
//
// -----------------------------------------------------------------------------
// File name:
// ----------
//
// tb_csd_add_subb.v
//
// -----------------------------------------------------------------------------
// History:
// --------
//
//    - 2016-04-16 - ilesser - Original version.
//
// -----------------------------------------------------------------------------

`define SIM_CLK_PERIOD_NS 10
`timescale 1ns/1ps

// *****************************************************************************
// Interface
// *****************************************************************************
module tb_csd_add_subb ();
// *****************************************************************************

// *****************************************************************************
// Architecture
// *****************************************************************************

   // -----------------------------------------------------
   // Testbench controlled variables and signals
   // -----------------------------------------------------
   localparam        W = 1;
   reg               tb_subb_a;
   reg               tb_subb_b;
   reg   [2*W-1:0]   tb_a;
   reg   [2*W-1:0]   tb_b;
   reg   [2*W-1:0]   tb_s;
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Testbecnch wiring
   // -----------------------------------------------------
   wire  [2*W-1:0]   wire_s;
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Transactors
   // -----------------------------------------------------
   // TODO: add bin2csd transactor
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Monitors
   // -----------------------------------------------------
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Checkers
   // -----------------------------------------------------
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Device under verifiacion
   // -----------------------------------------------------
   csd_add_subb #(
      .W(W)
   ) duv (
      .subb_a  (tb_subb_a),
      .subb_b  (tb_subb_b),
      .a       (tb_a),
      .b       (tb_b),
      .s       (wire_s)
   );
   // -----------------------------------------------------

// *****************************************************************************

endmodule

