// -----------------------------------------------------------------------------
//  Copyright (c) 2016 Microelectronics Lab. FIUBA.
//  All Rights Reserved.
//
//  The information contained in this file is confidential and proprietary.
//  Any reproduction, use or disclosure, in whole or in part, of this
//  program, including any attempt to obtain a human-readable version of this
//  program, without the express, prior written consent of Microelectronics Lab.
//  FIUBA is strictly prohibited.
//
// -----------------------------------------------------------------------------
// Description:
// ------------
//
// Testbech for bkm block.
//
// -----------------------------------------------------------------------------
// File name:
// ----------
//
// tb_bkm.v
//
// -----------------------------------------------------------------------------
// History:
// --------
//
//    - 2016-04-23 - ilesser - Original version.
//
// -----------------------------------------------------------------------------

`define SIM_CLK_PERIOD_NS 10
`timescale 1ns/1ps
`include "bkm_defs.vh"

// *****************************************************************************
// Interface
// *****************************************************************************
module tb_bkm ();
// *****************************************************************************

// *****************************************************************************
// Architecture
// *****************************************************************************

   // -----------------------------------------------------
   // Testbench controlled variables and signals
   // -----------------------------------------------------
   localparam        W     = 64;
   localparam        LOG2W = 6;
   localparam        N     = 64;
   localparam        LOG2N = 6;

   reg               tb_stop;
   reg               tb_clk;
   reg               tb_arst;
   reg               tb_srst;
   reg               tb_enable;

   reg               tb_start;
   reg               tb_mode;
   reg   [1:0]       tb_format;
   reg   [W-1:0]     tb_E_x;
   reg   [W-1:0]     tb_E_y;
   reg   [W-1:0]     tb_L_x;
   reg   [W-1:0]     tb_L_y;
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Testbecnch wiring
   // -----------------------------------------------------
   wire              bkm_done;
   wire  [`FSIZE-1:0]bkm_flags;
   wire  [W-1:0]     bkm_x;
   wire  [W-1:0]     bkm_y;
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Transactors
   // -----------------------------------------------------
   simlib_clk_osc #(
      // ----------------------------------------------
      // Parameters
      // ----------------------------------------------
      .CLK_PERIOD_NS(`SIM_CLK_PERIOD_NS)
   ) clk_osc (
      // ----------------------------------------------
      // Ports in
      // ----------------------------------------------
      .stop(tb_stop),
      // ----------------------------------------------
      // Ports out
      // ----------------------------------------------
      .clk_out(tb_clk)
   );
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Monitors
   // -----------------------------------------------------
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Checkers
   // -----------------------------------------------------
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Device under verifiacion
   // -----------------------------------------------------
   // -----------------------------------------------------
   // BKM Core
   // -----------------------------------------------------
   bkm #(
    // ----------------------------------
    // Parameters
    // ----------------------------------
      .W                   (W),
      .LOG2W               (LOG2W),
      .N                   (N),
      .LOG2N               (LOG2N)
   ) duv (
    // ----------------------------------
    // Clock, reset & enable inputs
    // ----------------------------------
      .clk                 (tb_clk),
      .arst                (tb_arst),
      .srst                (tb_srst),
      .enable              (tb_enable),
    // ----------------------------------
    // Data inputs
    // ----------------------------------
      .start               (tb_start),
      .mode                (tb_mode),
      .format              (tb_format),
      .E_x_in              (tb_E_x),
      .E_y_in              (tb_E_y),
      .L_x_in              (tb_L_x),
      .L_y_in              (tb_L_y),
    // ----------------------------------
    // Data outputs
    // ----------------------------------
      .X_out               (bkm_x),
      .Y_out               (bkm_y),
      .flags               (bkm_flags),
      .done                (bkm_done)
   );
   // -----------------------------------------------------

// *****************************************************************************

endmodule

