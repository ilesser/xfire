// -----------------------------------------------------------------------------
//  Copyright (c) 2016 Microelectronics Lab. FIUBA.
//  All Rights Reserved.
//
//  The information contained in this file is confidential and proprietary.
//  Any reproduction, use or disclosure, in whole or in part, of this
//  program, including any attempt to obtain a human-readable version of this
//  program, without the express, prior written consent of Microelectronics Lab.
//  FIUBA is strictly prohibited.
//
// -----------------------------------------------------------------------------
// Description:
// ------------
//
// Testbench for csd_add_subb block.
//
// -----------------------------------------------------------------------------
// File name:
// ----------
//
// tb_csd_add_subb.v
//
// -----------------------------------------------------------------------------
// History:
// --------
//
//    - 2016-04-16 - ilesser - Original version.
//
// -----------------------------------------------------------------------------

`define SIM_CLK_PERIOD_NS 10
`timescale 1ns/1ps

// *****************************************************************************
// Interface
// *****************************************************************************
module tb_csd_add_subb ();
// *****************************************************************************

// *****************************************************************************
// Architecture
// *****************************************************************************

   // -----------------------------------------------------
   // Testbench controlled variables and signals
   // -----------------------------------------------------
   localparam        W = 4;
   reg               tb_subb_x;
   reg               tb_subb_y;
   reg   [W-1:0]     tb_x_bin;
   reg   [W-1:0]     tb_y_bin;
   reg   [W-1:0]     tb_z_bin;
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Testbecnch wiring
   // -----------------------------------------------------
   wire              c_bin;
   wire  [W-1:0]     z_bin;
   wire  [2*W-1:0]   x_csd;
   wire  [2*W-1:0]   y_csd;
   wire  [1:0]       c_csd;
   wire  [2*W-1:0]   z_csd;
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Transactors
   // -----------------------------------------------------
   bin2csd #(
    // ----------------------------------
    // Parameters
    // ----------------------------------
      .W                   (W)
   ) bin2csd_x (
    // ----------------------------------
    // Data inputs
    // ----------------------------------
      .x                   (tb_x_bin),
    // ----------------------------------
    // Data outputs
    // ----------------------------------
      .y                   (x_csd)
   );

   bin2csd #(
    // ----------------------------------
    // Parameters
    // ----------------------------------
      .W                   (W)
   ) bin2csd_y (
    // ----------------------------------
    // Data inputs
    // ----------------------------------
      .x                   (tb_y_bin),
    // ----------------------------------
    // Data outputs
    // ----------------------------------
      .y                   (y_csd)
   );

   csd2bin #(
    // ----------------------------------
    // Parameters
    // ----------------------------------
      .W                   (W+1)
   ) csd2bin_z (
    // ----------------------------------
    // Data inputs
    // ----------------------------------
      .x                   ({c_csd, z_csd}),
    // ----------------------------------
    // Data outputs
    // ----------------------------------
      .y                   ({c_bin, z_bin})
   );

   // -----------------------------------------------------

   // -----------------------------------------------------
   // Monitors
   // -----------------------------------------------------
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Checkers
   // -----------------------------------------------------
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Device under verifiacion
   // -----------------------------------------------------
   csd_add_subb #(
      .W(W)
   ) duv (
      .subb_a  (tb_subb_x),
      .subb_b  (tb_subb_y),
      .a       (x_csd),
      .b       (y_csd),
      .c       (c_csd),
      .s       (z_csd)
   );
   // -----------------------------------------------------

// *****************************************************************************

endmodule

