// -----------------------------------------------------------------------------
//  Copyright (c) 2016 Microelectronics Lab. FIUBA.
//  All Rights Reserved.
//
//  The information contained in this file is confidential and proprietary.
//  Any reproduction, use or disclosure, in whole or in part, of this
//  program, including any attempt to obtain a human-readable version of this
//  program, without the express, prior written consent of Microelectronics Lab.
//  FIUBA is strictly prohibited.
//
// -----------------------------------------------------------------------------
// Description:
// ------------
//
// Barrel shifter testbench.
//
// -----------------------------------------------------------------------------
// File name:
// ----------
//
// tb_barrel_shifter.v
//
// -----------------------------------------------------------------------------
// History:
// --------
//
//    - 2016-04-25 - ilesser - Original version.
//
// -----------------------------------------------------------------------------

`define SIM_CLK_PERIOD_NS 10
`timescale 1ns/1ps

// *****************************************************************************
// Interface
// *****************************************************************************
module tb_barrel_shifter ();
// *****************************************************************************

// *****************************************************************************
// Architecture
// *****************************************************************************

   // -----------------------------------------------------
   // Testbench controlled variables and signals
   // -----------------------------------------------------
   localparam        W = 64;
   localparam        LOG2W = 6;
   reg               tb_dir;
   reg               tb_op;
   reg               tb_shift_t;
   reg   [LOG2W-1:0] tb_sel;
   reg   [W-1:0]     tb_in;
   reg   [W-1:0]     tb_out;
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Testbecnch wiring
   // -----------------------------------------------------
   wire  [W-1:0]     wire_out;
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Transactors
   // -----------------------------------------------------
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Monitors
   // -----------------------------------------------------
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Checkers
   // -----------------------------------------------------
   // -----------------------------------------------------

   // -----------------------------------------------------
   // Device under verifiacion
   // -----------------------------------------------------
   barrel_shifter #(
      .W(W),
      .LOG2W(LOG2W)
   ) duv (
      .dir(tb_dir),
      .op(tb_op),
      .shift_t(tb_shift_t),
      .in(tb_in),
      .out(wire_out)
   );
   // -----------------------------------------------------

// *****************************************************************************

endmodule

