//--------------------------------------------------------------------------------
//
// BKM LUT automatically generated on 11:23:34 AM (ART) Tuesday 13 September 2016
// using the bkm_lut.m function. Version = 1.2, from Saturday 08 September 2016.
// Parameters:
// Number of steps of the algorithm:            N     = 64
// Word size:                                   W     = 64
// Integer word size:                           WI    = 11
// Data channel upper guard bits:               UGD   = 2
// Integer word size of the data channel:       WDI   = 13
// Fractional word size of the data channel:    WDF   = 59
// Data channel lower guard bits:               LGD   = 6
// Word size of the data channel:               WD    = 72
// Control channel upper guard bits:            UGC   = 3
// Integer word size of the control channel:    WDI   = 14
// Fractional word size of the control channel: WDF   = 8
// Control channel lower guard bits:            LGC   = 4
// Word size of the control channel:            WC    = 22
//
//--------------------------------------------------------------------------------
//
//          IIIIIIIIIIIIIII.FFFFFFFFFFFFFF
//       +-----------------------------------+
// WD =  |  UGD   +  WI    +  W-WI  +  LGD   |
//       +-----------------------------------+
// WD =  |       WDI       +       WDF       |
//       +-----------------------------------+
//
//       +-----------------------------------+
// WC =  |  UGC   +   WI   +   4    +  LGC   |
//       +-----------------------------------+
// WC =  |       WCI       +       WCF       |
//       +-----------------------------------+
//          IIIIIIIIIIIIIII.FFFFFFFFFFFFFF
//
//--------------------------------------------------------------------------------
//
//
//--------------------------------------------------------------------------------
// This LUT uses 144 bits which represent 72 CSD digits. 
// They are represented by 36 hexadecimal digits. 
// After the LUT value you have the twos complement representation in 18 hexadecimal digits. 
// Since we use 13 bits for the integer part then the first 4.0 hexa digits represent the integer part. 
// The rest 14.0 hexa digits represent the fractional part.
// Example:
//sign X[4'bXXXX] [XX] = 144'h 040000000000000000000000000000000000;  // 200000000000000000 +1024.0000000000000000
//sign X[4'bXXXX] [XX] = 144'h 010000000000000000000000000000000000;  // 100000000000000000 +512.0000000000000000
//sign X[4'bXXXX] [XX] = 144'h 004000000000000000000000000000000000;  // 080000000000000000 +256.0000000000000000
//sign X[4'bXXXX] [XX] = 144'h 001000000000000000000000000000000000;  // 040000000000000000 +128.0000000000000000
//sign X[4'bXXXX] [XX] = 144'h 000400000000000000000000000000000000;  // 020000000000000000 +64.0000000000000000
//sign X[4'bXXXX] [XX] = 144'h 000100000000000000000000000000000000;  // 010000000000000000 +32.0000000000000000
//sign X[4'bXXXX] [XX] = 144'h 000040000000000000000000000000000000;  // 008000000000000000 +16.0000000000000000
//sign X[4'bXXXX] [XX] = 144'h 000010000000000000000000000000000000;  // 004000000000000000 +8.0000000000000000
//sign X[4'bXXXX] [XX] = 144'h 000004000000000000000000000000000000;  // 002000000000000000 +4.0000000000000000
//sign X[4'bXXXX] [XX] = 144'h 000001000000000000000000000000000000;  // 001000000000000000 +2.0000000000000000
//sign X[4'bXXXX] [XX] = 144'h 000000400000000000000000000000000000;  // 000800000000000000 +1.0000000000000000
//sign X[4'bXXXX] [XX] = 144'h 000000100000000000000000000000000000;  // 000400000000000000 +0.5000000000000000
//sign X[4'bXXXX] [XX] = 144'h 000000040000000000000000000000000000;  // 000200000000000000 +0.2500000000000000
//sign X[4'bXXXX] [XX] = 144'h 000000010000000000000000000000000000;  // 000100000000000000 +0.1250000000000000
//sign X[4'bXXXX] [XX] = 144'h 000000004000000000000000000000000000;  // 000080000000000000 +0.0625000000000000
//sign X[4'bXXXX] [XX] = 144'h 000000001000000000000000000000000000;  // 000040000000000000 +0.0312500000000000
//sign X[4'bXXXX] [XX] = 144'h 000000000400000000000000000000000000;  // 000020000000000000 +0.0156250000000000
//sign X[4'bXXXX] [XX] = 144'h 000000000100000000000000000000000000;  // 000010000000000000 +0.0078125000000000
//sign X[4'bXXXX] [XX] = 144'h 000000000040000000000000000000000000;  // 000008000000000000 +0.0039062500000000
//sign X[4'bXXXX] [XX] = 144'h 000000000010000000000000000000000000;  // 000004000000000000 +0.0019531250000000
//sign X[4'bXXXX] [XX] = 144'h 000000000004000000000000000000000000;  // 000002000000000000 +0.0009765625000000
//sign X[4'bXXXX] [XX] = 144'h 000000000001000000000000000000000000;  // 000001000000000000 +0.0004882812500000
//sign X[4'bXXXX] [XX] = 144'h 000000000000400000000000000000000000;  // 000000800000000000 +0.0002441406250000
//sign X[4'bXXXX] [XX] = 144'h 000000000000100000000000000000000000;  // 000000400000000000 +0.0001220703125000
//sign X[4'bXXXX] [XX] = 144'h 000000000000040000000000000000000000;  // 000000200000000000 +0.0000610351562500
//sign X[4'bXXXX] [XX] = 144'h 000000000000010000000000000000000000;  // 000000100000000000 +0.0000305175781250
//sign X[4'bXXXX] [XX] = 144'h 000000000000004000000000000000000000;  // 000000080000000000 +0.0000152587890625
//sign X[4'bXXXX] [XX] = 144'h 000000000000001000000000000000000000;  // 000000040000000000 +0.0000076293945312
//sign X[4'bXXXX] [XX] = 144'h 000000000000000400000000000000000000;  // 000000020000000000 +0.0000038146972656
//sign X[4'bXXXX] [XX] = 144'h 000000000000000100000000000000000000;  // 000000010000000000 +0.0000019073486328
//sign X[4'bXXXX] [XX] = 144'h 000000000000000040000000000000000000;  // 000000008000000000 +0.0000009536743164
//sign X[4'bXXXX] [XX] = 144'h 000000000000000010000000000000000000;  // 000000004000000000 +0.0000004768371582
//sign X[4'bXXXX] [XX] = 144'h 000000000000000004000000000000000000;  // 000000002000000000 +0.0000002384185791
//sign X[4'bXXXX] [XX] = 144'h 000000000000000001000000000000000000;  // 000000001000000000 +0.0000001192092896
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000400000000000000000;  // 000000000800000000 +0.0000000596046448
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000100000000000000000;  // 000000000400000000 +0.0000000298023224
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000040000000000000000;  // 000000000200000000 +0.0000000149011612
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000010000000000000000;  // 000000000100000000 +0.0000000074505806
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000004000000000000000;  // 000000000080000000 +0.0000000037252903
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000001000000000000000;  // 000000000040000000 +0.0000000018626451
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000400000000000000;  // 000000000020000000 +0.0000000009313226
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000100000000000000;  // 000000000010000000 +0.0000000004656613
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000040000000000000;  // 000000000008000000 +0.0000000002328306
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000010000000000000;  // 000000000004000000 +0.0000000001164153
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000004000000000000;  // 000000000002000000 +0.0000000000582077
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000001000000000000;  // 000000000001000000 +0.0000000000291038
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000400000000000;  // 000000000000800000 +0.0000000000145519
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000100000000000;  // 000000000000400000 +0.0000000000072760
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000040000000000;  // 000000000000200000 +0.0000000000036380
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000010000000000;  // 000000000000100000 +0.0000000000018190
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000004000000000;  // 000000000000080000 +0.0000000000009095
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000001000000000;  // 000000000000040000 +0.0000000000004547
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000000400000000;  // 000000000000020000 +0.0000000000002274
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000000100000000;  // 000000000000010000 +0.0000000000001137
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000000040000000;  // 000000000000008000 +0.0000000000000568
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000000010000000;  // 000000000000004000 +0.0000000000000284
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000000004000000;  // 000000000000002000 +0.0000000000000142
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000000001000000;  // 000000000000001000 +0.0000000000000071
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000000000400000;  // 000000000000000800 +0.0000000000000036
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000000000100000;  // 000000000000000400 +0.0000000000000018
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000000000040000;  // 000000000000000200 +0.0000000000000009
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000000000010000;  // 000000000000000100 +0.0000000000000004
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000000000004000;  // 000000000000000080 +0.0000000000000002
//sign X[4'bXXXX] [XX] = 144'h 000000000000000000000000000000001000;  // 000000000000000040 +0.0000000000000001
//--------------------------------------------------------------------------------
//
assign X[4'b0000] [01] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-1+1) + ( 0^2+ 0^2) * 2^(-2*1) )   n =  1   d_n = 0 
assign X[4'b0000] [02] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-2+1) + ( 0^2+ 0^2) * 2^(-2*2) )   n =  2   d_n = 0 
assign X[4'b0000] [03] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-3+1) + ( 0^2+ 0^2) * 2^(-2*3) )   n =  3   d_n = 0 
assign X[4'b0000] [04] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-4+1) + ( 0^2+ 0^2) * 2^(-2*4) )   n =  4   d_n = 0 
assign X[4'b0000] [05] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-5+1) + ( 0^2+ 0^2) * 2^(-2*5) )   n =  5   d_n = 0 
assign X[4'b0000] [06] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-6+1) + ( 0^2+ 0^2) * 2^(-2*6) )   n =  6   d_n = 0 
assign X[4'b0000] [07] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-7+1) + ( 0^2+ 0^2) * 2^(-2*7) )   n =  7   d_n = 0 
assign X[4'b0000] [08] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-8+1) + ( 0^2+ 0^2) * 2^(-2*8) )   n =  8   d_n = 0 
assign X[4'b0000] [09] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-9+1) + ( 0^2+ 0^2) * 2^(-2*9) )   n =  9   d_n = 0 
assign X[4'b0000] [10] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = 0 
assign X[4'b0000] [11] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = 0 
assign X[4'b0000] [12] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = 0 
assign X[4'b0000] [13] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = 0 
assign X[4'b0000] [14] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = 0 
assign X[4'b0000] [15] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = 0 
assign X[4'b0000] [16] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = 0 
assign X[4'b0000] [17] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = 0 
assign X[4'b0000] [18] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = 0 
assign X[4'b0000] [19] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = 0 
assign X[4'b0000] [20] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = 0 
assign X[4'b0000] [21] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = 0 
assign X[4'b0000] [22] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = 0 
assign X[4'b0000] [23] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = 0 
assign X[4'b0000] [24] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = 0 
assign X[4'b0000] [25] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = 0 
assign X[4'b0000] [26] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = 0 
assign X[4'b0000] [27] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = 0 
assign X[4'b0000] [28] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = 0 
assign X[4'b0000] [29] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = 0 
assign X[4'b0000] [30] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = 0 
assign X[4'b0000] [31] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = 0 
assign X[4'b0000] [32] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = 0 
assign X[4'b0000] [33] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = 0 
assign X[4'b0000] [34] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = 0 
assign X[4'b0000] [35] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = 0 
assign X[4'b0000] [36] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = 0 
assign X[4'b0000] [37] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = 0 
assign X[4'b0000] [38] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = 0 
assign X[4'b0000] [39] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = 0 
assign X[4'b0000] [40] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = 0 
assign X[4'b0000] [41] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = 0 
assign X[4'b0000] [42] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = 0 
assign X[4'b0000] [43] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = 0 
assign X[4'b0000] [44] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = 0 
assign X[4'b0000] [45] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = 0 
assign X[4'b0000] [46] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = 0 
assign X[4'b0000] [47] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = 0 
assign X[4'b0000] [48] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = 0 
assign X[4'b0000] [49] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = 0 
assign X[4'b0000] [50] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = 0 
assign X[4'b0000] [51] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = 0 
assign X[4'b0000] [52] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = 0 
assign X[4'b0000] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = 0 
assign X[4'b0000] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = 0 
assign X[4'b0000] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = 0 
assign X[4'b0000] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = 0 
assign X[4'b0000] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = 0 
assign X[4'b0000] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = 0 
assign X[4'b0000] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = 0 
assign X[4'b0000] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = 0 
assign X[4'b0000] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = 0 
assign X[4'b0000] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = 0 
assign X[4'b0000] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = 0 
assign X[4'b0000] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = 0 
assign X[4'b0001] [01] = 144'h 000000121008481040088480021200448000;  // 00033E647D97F30980 +0.4054651081081644 = 0.5 * ln( 1 +  1 * 2^(-1+1) + ( 1^2+ 0^2) * 2^(-2*1) )   n =  1   d_n = 1 
assign X[4'b0001] [02] = 144'h 000000042041000080204084844484040400;  // 0001C8FF7C79A9A220 +0.2231435513142098 = 0.5 * ln( 1 +  1 * 2^(-2+1) + ( 1^2+ 0^2) * 2^(-2*2) )   n =  2   d_n = 1 
assign X[4'b0001] [03] = 144'h 000000010201108010208204888084821200;  // 0000F1383B71579730 +0.1177830356563835 = 0.5 * ln( 1 +  1 * 2^(-3+1) + ( 1^2+ 0^2) * 2^(-2*3) )   n =  3   d_n = 1 
assign X[4'b0001] [04] = 144'h 000000004020044120120000104880444480;  // 00007C28C300458A98 +0.0606246218164348 = 0.5 * ln( 1 +  1 * 2^(-4+1) + ( 1^2+ 0^2) * 2^(-2*4) )   n =  4   d_n = 1 
assign X[4'b0001] [05] = 144'h 000000001002001110880421020048480000;  // 00003F05361CF06600 +0.0307716586667537 = 0.5 * ln( 1 +  1 * 2^(-5+1) + ( 1^2+ 0^2) * 2^(-2*5) )   n =  5   d_n = 1 
assign X[4'b0001] [06] = 144'h 000000000400200044412201002000100810;  // 00001FC0A8B0FC03E4 +0.0155041865359653 = 0.5 * ln( 1 +  1 * 2^(-6+1) + ( 1^2+ 0^2) * 2^(-2*6) )   n =  6   d_n = 1 
assign X[4'b0001] [07] = 144'h 000000000100020001111088804012102010;  // 00000FF015358833C4 +0.0077821404420549 = 0.5 * ln( 1 +  1 * 2^(-7+1) + ( 1^2+ 0^2) * 2^(-2*7) )   n =  7   d_n = 1 
assign X[4'b0001] [08] = 144'h 000000000040002000044441222010120200;  // 000007FC02A8AC42F0 +0.0038986404156573 = 0.5 * ln( 1 +  1 * 2^(-8+1) + ( 1^2+ 0^2) * 2^(-2*8) )   n =  8   d_n = 1 
assign X[4'b0001] [09] = 144'h 000000000010000200001111108888040421;  // 000003FF005535621C +0.0019512201312617 = 0.5 * ln( 1 +  1 * 2^(-9+1) + ( 1^2+ 0^2) * 2^(-2*9) )   n =  9   d_n = 1 
assign X[4'b0001] [10] = 144'h 000000000004000020000044444122220101;  // 000001FFC00AA8AB11 +0.0009760859730555 = 0.5 * ln( 1 +  1 * 2^(-10+1) + ( 1^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = 1 
assign X[4'b0001] [11] = 144'h 000000000001000002000001111110888880;  // 000000FFF001553558 +0.0004881620795014 = 0.5 * ln( 1 +  1 * 2^(-11+1) + ( 1^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = 1 
assign X[4'b0001] [12] = 144'h 000000000000400000200000044444412222;  // 0000007FFC002AA8AA +0.0002441108275274 = 0.5 * ln( 1 +  1 * 2^(-12+1) + ( 1^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = 1 
assign X[4'b0001] [13] = 144'h 000000000000100000020000001111111211;  // 0000003FFF00055535 +0.0001220628625257 = 0.5 * ln( 1 +  1 * 2^(-13+1) + ( 1^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = 1 
assign X[4'b0001] [14] = 144'h 000000000000040000002000000044444440;  // 0000001FFFC000AAA8 +0.0000610332936806 = 0.5 * ln( 1 +  1 * 2^(-14+1) + ( 1^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = 1 
assign X[4'b0001] [15] = 144'h 000000000000010000000200000001111111;  // 0000000FFFF0001555 +0.0000305171124732 = 0.5 * ln( 1 +  1 * 2^(-15+1) + ( 1^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = 1 
assign X[4'b0001] [16] = 144'h 000000000000004000000020000000044444;  // 00000007FFFC0002AA +0.0000152586726484 = 0.5 * ln( 1 +  1 * 2^(-16+1) + ( 1^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = 1 
assign X[4'b0001] [17] = 144'h 000000000000001000000002000000001111;  // 00000003FFFF000055 +0.0000076293654276 = 0.5 * ln( 1 +  1 * 2^(-17+1) + ( 1^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = 1 
assign X[4'b0001] [18] = 144'h 000000000000000400000000200000000044;  // 00000001FFFFC0000A +0.0000038146899897 = 0.5 * ln( 1 +  1 * 2^(-18+1) + ( 1^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = 1 
assign X[4'b0001] [19] = 144'h 000000000000000100000000020000000001;  // 00000000FFFFF00001 +0.0000019073468138 = 0.5 * ln( 1 +  1 * 2^(-19+1) + ( 1^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = 1 
assign X[4'b0001] [20] = 144'h 000000000000000040000000002000000000;  // 000000007FFFFC0000 +0.0000009536738617 = 0.5 * ln( 1 +  1 * 2^(-20+1) + ( 1^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = 1 
assign X[4'b0001] [21] = 144'h 000000000000000010000000000200000000;  // 000000003FFFFF0000 +0.0000004768370445 = 0.5 * ln( 1 +  1 * 2^(-21+1) + ( 1^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = 1 
assign X[4'b0001] [22] = 144'h 000000000000000004000000000020000000;  // 000000001FFFFFC000 +0.0000002384185507 = 0.5 * ln( 1 +  1 * 2^(-22+1) + ( 1^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = 1 
assign X[4'b0001] [23] = 144'h 000000000000000001000000000002000000;  // 000000000FFFFFF000 +0.0000001192092824 = 0.5 * ln( 1 +  1 * 2^(-23+1) + ( 1^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = 1 
assign X[4'b0001] [24] = 144'h 000000000000000000400000000000200000;  // 0000000007FFFFFC00 +0.0000000596046430 = 0.5 * ln( 1 +  1 * 2^(-24+1) + ( 1^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = 1 
assign X[4'b0001] [25] = 144'h 000000000000000000100000000000020000;  // 0000000003FFFFFF00 +0.0000000298023219 = 0.5 * ln( 1 +  1 * 2^(-25+1) + ( 1^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = 1 
assign X[4'b0001] [26] = 144'h 000000000000000000040000000000002000;  // 0000000001FFFFFFC0 +0.0000000149011611 = 0.5 * ln( 1 +  1 * 2^(-26+1) + ( 1^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = 1 
assign X[4'b0001] [27] = 144'h 000000000000000000010000000000000200;  // 0000000000FFFFFFF0 +0.0000000074505806 = 0.5 * ln( 1 +  1 * 2^(-27+1) + ( 1^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = 1 
assign X[4'b0001] [28] = 144'h 000000000000000000004000000000000020;  // 00000000007FFFFFFC +0.0000000037252903 = 0.5 * ln( 1 +  1 * 2^(-28+1) + ( 1^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = 1 
assign X[4'b0001] [29] = 144'h 000000000000000000001000000000000002;  // 00000000003FFFFFFF +0.0000000018626451 = 0.5 * ln( 1 +  1 * 2^(-29+1) + ( 1^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = 1 
assign X[4'b0001] [30] = 144'h 000000000000000000000400000000000000;  // 00000000001FFFFFFF +0.0000000009313226 = 0.5 * ln( 1 +  1 * 2^(-30+1) + ( 1^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = 1 
assign X[4'b0001] [31] = 144'h 000000000000000000000100000000000000;  // 00000000000FFFFFFF +0.0000000004656613 = 0.5 * ln( 1 +  1 * 2^(-31+1) + ( 1^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = 1 
assign X[4'b0001] [32] = 144'h 000000000000000000000040000000000000;  // 000000000007FFFFFF +0.0000000002328306 = 0.5 * ln( 1 +  1 * 2^(-32+1) + ( 1^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = 1 
assign X[4'b0001] [33] = 144'h 000000000000000000000010000000000000;  // 000000000003FFFFFF +0.0000000001164153 = 0.5 * ln( 1 +  1 * 2^(-33+1) + ( 1^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = 1 
assign X[4'b0001] [34] = 144'h 000000000000000000000004000000000000;  // 000000000001FFFFFF +0.0000000000582077 = 0.5 * ln( 1 +  1 * 2^(-34+1) + ( 1^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = 1 
assign X[4'b0001] [35] = 144'h 000000000000000000000001000000000000;  // 000000000000FFFFFF +0.0000000000291038 = 0.5 * ln( 1 +  1 * 2^(-35+1) + ( 1^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = 1 
assign X[4'b0001] [36] = 144'h 000000000000000000000000400000000000;  // 0000000000007FFFFF +0.0000000000145519 = 0.5 * ln( 1 +  1 * 2^(-36+1) + ( 1^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = 1 
assign X[4'b0001] [37] = 144'h 000000000000000000000000100000000000;  // 0000000000003FFFFF +0.0000000000072760 = 0.5 * ln( 1 +  1 * 2^(-37+1) + ( 1^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = 1 
assign X[4'b0001] [38] = 144'h 000000000000000000000000040000000000;  // 0000000000001FFFFF +0.0000000000036380 = 0.5 * ln( 1 +  1 * 2^(-38+1) + ( 1^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = 1 
assign X[4'b0001] [39] = 144'h 000000000000000000000000010000000000;  // 0000000000000FFFFF +0.0000000000018190 = 0.5 * ln( 1 +  1 * 2^(-39+1) + ( 1^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = 1 
assign X[4'b0001] [40] = 144'h 000000000000000000000000004000000000;  // 00000000000007FFFF +0.0000000000009095 = 0.5 * ln( 1 +  1 * 2^(-40+1) + ( 1^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = 1 
assign X[4'b0001] [41] = 144'h 000000000000000000000000001000000000;  // 00000000000003FFFF +0.0000000000004547 = 0.5 * ln( 1 +  1 * 2^(-41+1) + ( 1^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = 1 
assign X[4'b0001] [42] = 144'h 000000000000000000000000000400000000;  // 00000000000001FFFF +0.0000000000002274 = 0.5 * ln( 1 +  1 * 2^(-42+1) + ( 1^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = 1 
assign X[4'b0001] [43] = 144'h 000000000000000000000000000100000000;  // 00000000000000FFFF +0.0000000000001137 = 0.5 * ln( 1 +  1 * 2^(-43+1) + ( 1^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = 1 
assign X[4'b0001] [44] = 144'h 000000000000000000000000000040000000;  // 000000000000007FFF +0.0000000000000568 = 0.5 * ln( 1 +  1 * 2^(-44+1) + ( 1^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = 1 
assign X[4'b0001] [45] = 144'h 000000000000000000000000000010000000;  // 000000000000003FFF +0.0000000000000284 = 0.5 * ln( 1 +  1 * 2^(-45+1) + ( 1^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = 1 
assign X[4'b0001] [46] = 144'h 000000000000000000000000000004000000;  // 000000000000001FFF +0.0000000000000142 = 0.5 * ln( 1 +  1 * 2^(-46+1) + ( 1^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = 1 
assign X[4'b0001] [47] = 144'h 000000000000000000000000000001000000;  // 000000000000000FFF +0.0000000000000071 = 0.5 * ln( 1 +  1 * 2^(-47+1) + ( 1^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = 1 
assign X[4'b0001] [48] = 144'h 000000000000000000000000000000400000;  // 0000000000000007FF +0.0000000000000036 = 0.5 * ln( 1 +  1 * 2^(-48+1) + ( 1^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = 1 
assign X[4'b0001] [49] = 144'h 000000000000000000000000000000100000;  // 0000000000000003FF +0.0000000000000018 = 0.5 * ln( 1 +  1 * 2^(-49+1) + ( 1^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = 1 
assign X[4'b0001] [50] = 144'h 000000000000000000000000000000040000;  // 0000000000000001FF +0.0000000000000009 = 0.5 * ln( 1 +  1 * 2^(-50+1) + ( 1^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = 1 
assign X[4'b0001] [51] = 144'h 000000000000000000000000000000010000;  // 0000000000000000FF +0.0000000000000004 = 0.5 * ln( 1 +  1 * 2^(-51+1) + ( 1^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = 1 
assign X[4'b0001] [52] = 144'h 000000000000000000000000000000004000;  // 00000000000000007F +0.0000000000000002 = 0.5 * ln( 1 +  1 * 2^(-52+1) + ( 1^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = 1 
assign X[4'b0001] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-53+1) + ( 1^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = 1 
assign X[4'b0001] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-54+1) + ( 1^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = 1 
assign X[4'b0001] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-55+1) + ( 1^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = 1 
assign X[4'b0001] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-56+1) + ( 1^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = 1 
assign X[4'b0001] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-57+1) + ( 1^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = 1 
assign X[4'b0001] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-58+1) + ( 1^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = 1 
assign X[4'b0001] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-59+1) + ( 1^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = 1 
assign X[4'b0001] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-60+1) + ( 1^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = 1 
assign X[4'b0001] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-61+1) + ( 1^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = 1 
assign X[4'b0001] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-62+1) + ( 1^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = 1 
assign X[4'b0001] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-63+1) + ( 1^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = 1 
assign X[4'b0001] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-64+1) + ( 1^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = 1 
assign X[4'b0010] [01] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-1+1) + ( 0^2+ 0^2) * 2^(-2*1) )   n =  1   d_n = -0 
assign X[4'b0010] [02] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-2+1) + ( 0^2+ 0^2) * 2^(-2*2) )   n =  2   d_n = -0 
assign X[4'b0010] [03] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-3+1) + ( 0^2+ 0^2) * 2^(-2*3) )   n =  3   d_n = -0 
assign X[4'b0010] [04] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-4+1) + ( 0^2+ 0^2) * 2^(-2*4) )   n =  4   d_n = -0 
assign X[4'b0010] [05] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-5+1) + ( 0^2+ 0^2) * 2^(-2*5) )   n =  5   d_n = -0 
assign X[4'b0010] [06] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-6+1) + ( 0^2+ 0^2) * 2^(-2*6) )   n =  6   d_n = -0 
assign X[4'b0010] [07] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-7+1) + ( 0^2+ 0^2) * 2^(-2*7) )   n =  7   d_n = -0 
assign X[4'b0010] [08] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-8+1) + ( 0^2+ 0^2) * 2^(-2*8) )   n =  8   d_n = -0 
assign X[4'b0010] [09] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-9+1) + ( 0^2+ 0^2) * 2^(-2*9) )   n =  9   d_n = -0 
assign X[4'b0010] [10] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = -0 
assign X[4'b0010] [11] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = -0 
assign X[4'b0010] [12] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = -0 
assign X[4'b0010] [13] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = -0 
assign X[4'b0010] [14] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = -0 
assign X[4'b0010] [15] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = -0 
assign X[4'b0010] [16] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = -0 
assign X[4'b0010] [17] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = -0 
assign X[4'b0010] [18] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = -0 
assign X[4'b0010] [19] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = -0 
assign X[4'b0010] [20] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = -0 
assign X[4'b0010] [21] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = -0 
assign X[4'b0010] [22] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = -0 
assign X[4'b0010] [23] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = -0 
assign X[4'b0010] [24] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = -0 
assign X[4'b0010] [25] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = -0 
assign X[4'b0010] [26] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = -0 
assign X[4'b0010] [27] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = -0 
assign X[4'b0010] [28] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = -0 
assign X[4'b0010] [29] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = -0 
assign X[4'b0010] [30] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = -0 
assign X[4'b0010] [31] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = -0 
assign X[4'b0010] [32] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = -0 
assign X[4'b0010] [33] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = -0 
assign X[4'b0010] [34] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = -0 
assign X[4'b0010] [35] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = -0 
assign X[4'b0010] [36] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = -0 
assign X[4'b0010] [37] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = -0 
assign X[4'b0010] [38] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = -0 
assign X[4'b0010] [39] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = -0 
assign X[4'b0010] [40] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = -0 
assign X[4'b0010] [41] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = -0 
assign X[4'b0010] [42] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = -0 
assign X[4'b0010] [43] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = -0 
assign X[4'b0010] [44] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = -0 
assign X[4'b0010] [45] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = -0 
assign X[4'b0010] [46] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = -0 
assign X[4'b0010] [47] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = -0 
assign X[4'b0010] [48] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = -0 
assign X[4'b0010] [49] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = -0 
assign X[4'b0010] [50] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = -0 
assign X[4'b0010] [51] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = -0 
assign X[4'b0010] [52] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = -0 
assign X[4'b0010] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = -0 
assign X[4'b0010] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = -0 
assign X[4'b0010] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = -0 
assign X[4'b0010] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = -0 
assign X[4'b0010] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = -0 
assign X[4'b0010] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = -0 
assign X[4'b0010] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = -0 
assign X[4'b0010] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = -0 
assign X[4'b0010] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = -0 
assign X[4'b0010] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = -0 
assign X[4'b0010] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = -0 
assign X[4'b0010] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = -0 
assign X[4'b0011] [01] = 144'h 000000844210420210001004820480101000;  // FFFA746F4041700000 -0.6931471805599453 = 0.5 * ln( 1 + -1 * 2^(-1+1) + (-1^2+ 0^2) * 2^(-2*1) )   n =  1   d_n = -1 
assign X[4'b0011] [02] = 144'h 000000082212211020080884881041082000;  // FFFDB2D3BDD9680000 -0.2876820724517809 = 0.5 * ln( 1 + -1 * 2^(-2+1) + (-1^2+ 0^2) * 2^(-2*2) )   n =  2   d_n = -1 
assign X[4'b0011] [03] = 144'h 000000020208404204800808800420801000;  // FFFEEE8717DD800000 -0.1335313926245226 = 0.5 * ln( 1 + -1 * 2^(-3+1) + (-1^2+ 0^2) * 2^(-2*3) )   n =  3   d_n = -1 
assign X[4'b0011] [04] = 144'h 000000008020211210841112010812002040;  // FFFF7BD33A53100000 -0.0645385211375712 = 0.5 * ln( 1 + -1 * 2^(-4+1) + (-1^2+ 0^2) * 2^(-2*4) )   n =  4   d_n = -1 
assign X[4'b0011] [05] = 144'h 000000002002008440440880481202020200;  // FFFFBEFA89D8600000 -0.0317486983145803 = 0.5 * ln( 1 + -1 * 2^(-5+1) + (-1^2+ 0^2) * 2^(-2*5) )   n =  5   d_n = -1 
assign X[4'b0011] [06] = 144'h 000000000800200211121102088111008204;  // FFFFDFBF534ED80000 -0.0157483569681392 = 0.5 * ln( 1 + -1 * 2^(-6+1) + (-1^2+ 0^2) * 2^(-2*6) )   n =  6   d_n = -1 
assign X[4'b0011] [07] = 144'h 000000000200020008444044408204048102;  // FFFFEFEFEA8A780000 -0.0078431774610259 = 0.5 * ln( 1 + -1 * 2^(-7+1) + (-1^2+ 0^2) * 2^(-2*7) )   n =  7   d_n = -1 
assign X[4'b0011] [08] = 144'h 000000000080002000211112111020844848;  // FFFFF7FBFD53500000 -0.0039138993211363 = 0.5 * ln( 1 + -1 * 2^(-8+1) + (-1^2+ 0^2) * 2^(-2*8) )   n =  8   d_n = -1 
assign X[4'b0011] [09] = 144'h 000000000020000200008444404444080880;  // FFFFFBFEFFAA880000 -0.0019550348358034 = 0.5 * ln( 1 + -1 * 2^(-9+1) + (-1^2+ 0^2) * 2^(-2*9) )   n =  9   d_n = -1 
assign X[4'b0011] [10] = 144'h 000000000008000020000211111211110202;  // FFFFFDFFBFF5500000 -0.0009770396478266 = 0.5 * ln( 1 + -1 * 2^(-10+1) + (-1^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = -1 
assign X[4'b0011] [11] = 144'h 000000000002000002000008444440444440;  // FFFFFEFFEFFEA80000 -0.0004884004981089 = 0.5 * ln( 1 + -1 * 2^(-11+1) + (-1^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = -1 
assign X[4'b0011] [12] = 144'h 000000000000800000200000211111121111;  // FFFFFF7FFBFFD80000 -0.0002441704321739 = 0.5 * ln( 1 + -1 * 2^(-12+1) + (-1^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = -1 
assign X[4'b0011] [13] = 144'h 000000000000200000020000008444444044;  // FFFFFFBFFEFFF80000 -0.0001220777636870 = 0.5 * ln( 1 + -1 * 2^(-13+1) + (-1^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = -1 
assign X[4'b0011] [14] = 144'h 000000000000080000002000000211111110;  // FFFFFFDFFFC0000000 -0.0000610370189709 = 0.5 * ln( 1 + -1 * 2^(-14+1) + (-1^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = -1 
assign X[4'b0011] [15] = 144'h 000000000000020000000200000008444444;  // FFFFFFEFFFF0000000 -0.0000305180437958 = 0.5 * ln( 1 + -1 * 2^(-15+1) + (-1^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = -1 
assign X[4'b0011] [16] = 144'h 000000000000008000000020000000088888;  // FFFFFFF7FFFC000000 -0.0000152589054790 = 0.5 * ln( 1 + -1 * 2^(-16+1) + (-1^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = -1 
assign X[4'b0011] [17] = 144'h 000000000000002000000002000000002222;  // FFFFFFFBFFFF000000 -0.0000076294236352 = 0.5 * ln( 1 + -1 * 2^(-17+1) + (-1^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = -1 
assign X[4'b0011] [18] = 144'h 000000000000000800000000200000000088;  // FFFFFFFDFFFFC00000 -0.0000038147045416 = 0.5 * ln( 1 + -1 * 2^(-18+1) + (-1^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = -1 
assign X[4'b0011] [19] = 144'h 000000000000000200000000020000000002;  // FFFFFFFEFFFFF00000 -0.0000019073504518 = 0.5 * ln( 1 + -1 * 2^(-19+1) + (-1^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = -1 
assign X[4'b0011] [20] = 144'h 000000000000000080000000002000000000;  // FFFFFFFF7FFFF80000 -0.0000009536747712 = 0.5 * ln( 1 + -1 * 2^(-20+1) + (-1^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = -1 
assign X[4'b0011] [21] = 144'h 000000000000000020000000000200000000;  // FFFFFFFFC000000000 -0.0000004768372719 = 0.5 * ln( 1 + -1 * 2^(-21+1) + (-1^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = -1 
assign X[4'b0011] [22] = 144'h 000000000000000008000000000020000000;  // FFFFFFFFE000000000 -0.0000002384186075 = 0.5 * ln( 1 + -1 * 2^(-22+1) + (-1^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = -1 
assign X[4'b0011] [23] = 144'h 000000000000000002000000000002000000;  // FFFFFFFFF000000000 -0.0000001192092967 = 0.5 * ln( 1 + -1 * 2^(-23+1) + (-1^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = -1 
assign X[4'b0011] [24] = 144'h 000000000000000000800000000000200000;  // FFFFFFFFF800000000 -0.0000000596046466 = 0.5 * ln( 1 + -1 * 2^(-24+1) + (-1^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = -1 
assign X[4'b0011] [25] = 144'h 000000000000000000200000000000020000;  // FFFFFFFFFC00000000 -0.0000000298023228 = 0.5 * ln( 1 + -1 * 2^(-25+1) + (-1^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = -1 
assign X[4'b0011] [26] = 144'h 000000000000000000080000000000002000;  // FFFFFFFFFE00000000 -0.0000000149011613 = 0.5 * ln( 1 + -1 * 2^(-26+1) + (-1^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = -1 
assign X[4'b0011] [27] = 144'h 000000000000000000020000000000000200;  // FFFFFFFFFF00000000 -0.0000000074505806 = 0.5 * ln( 1 + -1 * 2^(-27+1) + (-1^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = -1 
assign X[4'b0011] [28] = 144'h 000000000000000000008000000000000020;  // FFFFFFFFFF80000000 -0.0000000037252903 = 0.5 * ln( 1 + -1 * 2^(-28+1) + (-1^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = -1 
assign X[4'b0011] [29] = 144'h 000000000000000000002000000000000002;  // FFFFFFFFFFC0000000 -0.0000000018626452 = 0.5 * ln( 1 + -1 * 2^(-29+1) + (-1^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = -1 
assign X[4'b0011] [30] = 144'h 000000000000000000000800000000000000;  // FFFFFFFFFFE0000000 -0.0000000009313226 = 0.5 * ln( 1 + -1 * 2^(-30+1) + (-1^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = -1 
assign X[4'b0011] [31] = 144'h 000000000000000000000200000000000000;  // FFFFFFFFFFF0000000 -0.0000000004656613 = 0.5 * ln( 1 + -1 * 2^(-31+1) + (-1^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = -1 
assign X[4'b0011] [32] = 144'h 000000000000000000000080000000000000;  // FFFFFFFFFFF8000000 -0.0000000002328306 = 0.5 * ln( 1 + -1 * 2^(-32+1) + (-1^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = -1 
assign X[4'b0011] [33] = 144'h 000000000000000000000020000000000000;  // FFFFFFFFFFFC000000 -0.0000000001164153 = 0.5 * ln( 1 + -1 * 2^(-33+1) + (-1^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = -1 
assign X[4'b0011] [34] = 144'h 000000000000000000000008000000000000;  // FFFFFFFFFFFE000000 -0.0000000000582077 = 0.5 * ln( 1 + -1 * 2^(-34+1) + (-1^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = -1 
assign X[4'b0011] [35] = 144'h 000000000000000000000002000000000000;  // FFFFFFFFFFFF000000 -0.0000000000291038 = 0.5 * ln( 1 + -1 * 2^(-35+1) + (-1^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = -1 
assign X[4'b0011] [36] = 144'h 000000000000000000000000800000000000;  // FFFFFFFFFFFF800000 -0.0000000000145519 = 0.5 * ln( 1 + -1 * 2^(-36+1) + (-1^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = -1 
assign X[4'b0011] [37] = 144'h 000000000000000000000000200000000000;  // FFFFFFFFFFFFC00000 -0.0000000000072760 = 0.5 * ln( 1 + -1 * 2^(-37+1) + (-1^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = -1 
assign X[4'b0011] [38] = 144'h 000000000000000000000000080000000000;  // FFFFFFFFFFFFE00000 -0.0000000000036380 = 0.5 * ln( 1 + -1 * 2^(-38+1) + (-1^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = -1 
assign X[4'b0011] [39] = 144'h 000000000000000000000000020000000000;  // FFFFFFFFFFFFF00000 -0.0000000000018190 = 0.5 * ln( 1 + -1 * 2^(-39+1) + (-1^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = -1 
assign X[4'b0011] [40] = 144'h 000000000000000000000000008000000000;  // FFFFFFFFFFFFF80000 -0.0000000000009095 = 0.5 * ln( 1 + -1 * 2^(-40+1) + (-1^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = -1 
assign X[4'b0011] [41] = 144'h 000000000000000000000000002000000000;  // FFFFFFFFFFFFF80000 -0.0000000000004547 = 0.5 * ln( 1 + -1 * 2^(-41+1) + (-1^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = -1 
assign X[4'b0011] [42] = 144'h 000000000000000000000000000800000000;  // 1000000000000000000 -0.0000000000002274 = 0.5 * ln( 1 + -1 * 2^(-42+1) + (-1^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = -1 
assign X[4'b0011] [43] = 144'h 000000000000000000000000000200000000;  // 1000000000000000000 -0.0000000000001137 = 0.5 * ln( 1 + -1 * 2^(-43+1) + (-1^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = -1 
assign X[4'b0011] [44] = 144'h 000000000000000000000000000080000000;  // 1000000000000000000 -0.0000000000000568 = 0.5 * ln( 1 + -1 * 2^(-44+1) + (-1^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = -1 
assign X[4'b0011] [45] = 144'h 000000000000000000000000000020000000;  // 1000000000000000000 -0.0000000000000284 = 0.5 * ln( 1 + -1 * 2^(-45+1) + (-1^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = -1 
assign X[4'b0011] [46] = 144'h 000000000000000000000000000008000000;  // 1000000000000000000 -0.0000000000000142 = 0.5 * ln( 1 + -1 * 2^(-46+1) + (-1^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = -1 
assign X[4'b0011] [47] = 144'h 000000000000000000000000000002000000;  // 1000000000000000000 -0.0000000000000071 = 0.5 * ln( 1 + -1 * 2^(-47+1) + (-1^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = -1 
assign X[4'b0011] [48] = 144'h 000000000000000000000000000000800000;  // 1000000000000000000 -0.0000000000000036 = 0.5 * ln( 1 + -1 * 2^(-48+1) + (-1^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = -1 
assign X[4'b0011] [49] = 144'h 000000000000000000000000000000200000;  // 1000000000000000000 -0.0000000000000018 = 0.5 * ln( 1 + -1 * 2^(-49+1) + (-1^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = -1 
assign X[4'b0011] [50] = 144'h 000000000000000000000000000000080000;  // 1000000000000000000 -0.0000000000000009 = 0.5 * ln( 1 + -1 * 2^(-50+1) + (-1^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = -1 
assign X[4'b0011] [51] = 144'h 000000000000000000000000000000020000;  // 1000000000000000000 -0.0000000000000004 = 0.5 * ln( 1 + -1 * 2^(-51+1) + (-1^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = -1 
assign X[4'b0011] [52] = 144'h 000000000000000000000000000000008000;  // 1000000000000000000 -0.0000000000000002 = 0.5 * ln( 1 + -1 * 2^(-52+1) + (-1^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = -1 
assign X[4'b0011] [53] = 144'h 000000000000000000000000000000002000;  // 1000000000000000000 -0.0000000000000001 = 0.5 * ln( 1 + -1 * 2^(-53+1) + (-1^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = -1 
assign X[4'b0011] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-54+1) + (-1^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = -1 
assign X[4'b0011] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-55+1) + (-1^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = -1 
assign X[4'b0011] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-56+1) + (-1^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = -1 
assign X[4'b0011] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-57+1) + (-1^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = -1 
assign X[4'b0011] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-58+1) + (-1^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = -1 
assign X[4'b0011] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-59+1) + (-1^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = -1 
assign X[4'b0011] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-60+1) + (-1^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = -1 
assign X[4'b0011] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-61+1) + (-1^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = -1 
assign X[4'b0011] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-62+1) + (-1^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = -1 
assign X[4'b0011] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-63+1) + (-1^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = -1 
assign X[4'b0011] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-64+1) + (-1^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = -1 
assign X[4'b0100] [01] = 144'h 000000010810400020081021211121010400;  // 0000E47FBE3CD4D128 +0.1115717756571049 = 0.5 * ln( 1 +  0 * 2^(-1+1) + ( 0^2+ 1^2) * 2^(-2*1) )   n =  1   d_n = 0+1i 
assign X[4'b0100] [02] = 144'h 000000001008011048048000041220111100;  // 00003E14618022C552 +0.0303123109082174 = 0.5 * ln( 1 +  0 * 2^(-2+1) + ( 0^2+ 1^2) * 2^(-2*2) )   n =  2   d_n = 0+1i 
assign X[4'b0100] [03] = 144'h 000000000100080011104880400800042120;  // 00000FE054587E01CC +0.0077520932679826 = 0.5 * ln( 1 +  0 * 2^(-3+1) + ( 0^2+ 1^2) * 2^(-2*3) )   n =  3   d_n = 0+1i 
assign X[4'b0100] [04] = 144'h 000000000010000800011110488804048404;  // 000003FE01545621A1 +0.0019493202078287 = 0.5 * ln( 1 +  0 * 2^(-4+1) + ( 0^2+ 1^2) * 2^(-2*4) )   n =  4   d_n = 0+1i 
assign X[4'b0100] [05] = 144'h 000000000001000008000011111048888084;  // 000000FFE00554557A +0.0004880429865277 = 0.5 * ln( 1 +  0 * 2^(-5+1) + ( 0^2+ 1^2) * 2^(-2*5) )   n =  5   d_n = 0+1i 
assign X[4'b0100] [06] = 144'h 000000000000100000080000011111100448;  // 0000003FFE00155425 +0.0001220554137636 = 0.5 * ln( 1 +  0 * 2^(-6+1) + ( 0^2+ 1^2) * 2^(-2*6) )   n =  6   d_n = 0+1i 
assign X[4'b0100] [07] = 144'h 000000000000010000000800000011111110;  // 0000000FFFE0005554 +0.0000305166468403 = 0.5 * ln( 1 +  0 * 2^(-7+1) + ( 0^2+ 1^2) * 2^(-2*7) )   n =  7   d_n = 0+1i 
assign X[4'b0100] [08] = 144'h 000000000000001000000008000000011111;  // 00000003FFFE000155 +0.0000076293363242 = 0.5 * ln( 1 +  0 * 2^(-8+1) + ( 0^2+ 1^2) * 2^(-2*8) )   n =  8   d_n = 0+1i 
assign X[4'b0100] [09] = 144'h 000000000000000100000000080000000012;  // 00000000FFFFE00003 +0.0000019073449948 = 0.5 * ln( 1 +  0 * 2^(-9+1) + ( 0^2+ 1^2) * 2^(-2*9) )   n =  9   d_n = 0+1i 
assign X[4'b0100] [10] = 144'h 000000000000000010000000000800000000;  // 000000003FFFFE0000 +0.0000004768369308 = 0.5 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 1^2) * 2^(-2*10) )   n = 10   d_n = 0+1i 
assign X[4'b0100] [11] = 144'h 000000000000000001000000000008000000;  // 000000000FFFFFE000 +0.0000001192092753 = 0.5 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 1^2) * 2^(-2*11) )   n = 11   d_n = 0+1i 
assign X[4'b0100] [12] = 144'h 000000000000000000100000000000080000;  // 0000000003FFFFFE00 +0.0000000298023215 = 0.5 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 1^2) * 2^(-2*12) )   n = 12   d_n = 0+1i 
assign X[4'b0100] [13] = 144'h 000000000000000000010000000000000200;  // 0000000000FFFFFFF0 +0.0000000074505806 = 0.5 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 1^2) * 2^(-2*13) )   n = 13   d_n = 0+1i 
assign X[4'b0100] [14] = 144'h 000000000000000000001000000000000002;  // 00000000003FFFFFFF +0.0000000018626451 = 0.5 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 1^2) * 2^(-2*14) )   n = 14   d_n = 0+1i 
assign X[4'b0100] [15] = 144'h 000000000000000000000100000000000000;  // 00000000000FFFFFFF +0.0000000004656613 = 0.5 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 1^2) * 2^(-2*15) )   n = 15   d_n = 0+1i 
assign X[4'b0100] [16] = 144'h 000000000000000000000010000000000000;  // 000000000003FFFFFF +0.0000000001164153 = 0.5 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 1^2) * 2^(-2*16) )   n = 16   d_n = 0+1i 
assign X[4'b0100] [17] = 144'h 000000000000000000000001000000000000;  // 000000000000FFFFFF +0.0000000000291038 = 0.5 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 1^2) * 2^(-2*17) )   n = 17   d_n = 0+1i 
assign X[4'b0100] [18] = 144'h 000000000000000000000000100000000000;  // 0000000000003FFFFF +0.0000000000072760 = 0.5 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 1^2) * 2^(-2*18) )   n = 18   d_n = 0+1i 
assign X[4'b0100] [19] = 144'h 000000000000000000000000010000000000;  // 0000000000000FFFFF +0.0000000000018190 = 0.5 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 1^2) * 2^(-2*19) )   n = 19   d_n = 0+1i 
assign X[4'b0100] [20] = 144'h 000000000000000000000000001000000000;  // 00000000000003FFFF +0.0000000000004547 = 0.5 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 1^2) * 2^(-2*20) )   n = 20   d_n = 0+1i 
assign X[4'b0100] [21] = 144'h 000000000000000000000000000100000000;  // 00000000000000FFFF +0.0000000000001137 = 0.5 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 1^2) * 2^(-2*21) )   n = 21   d_n = 0+1i 
assign X[4'b0100] [22] = 144'h 000000000000000000000000000010000000;  // 000000000000003FFF +0.0000000000000284 = 0.5 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 1^2) * 2^(-2*22) )   n = 22   d_n = 0+1i 
assign X[4'b0100] [23] = 144'h 000000000000000000000000000001000000;  // 000000000000000FFF +0.0000000000000071 = 0.5 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 1^2) * 2^(-2*23) )   n = 23   d_n = 0+1i 
assign X[4'b0100] [24] = 144'h 000000000000000000000000000000100000;  // 0000000000000003FF +0.0000000000000018 = 0.5 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 1^2) * 2^(-2*24) )   n = 24   d_n = 0+1i 
assign X[4'b0100] [25] = 144'h 000000000000000000000000000000010000;  // 0000000000000000FF +0.0000000000000004 = 0.5 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 1^2) * 2^(-2*25) )   n = 25   d_n = 0+1i 
assign X[4'b0100] [26] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 1^2) * 2^(-2*26) )   n = 26   d_n = 0+1i 
assign X[4'b0100] [27] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 1^2) * 2^(-2*27) )   n = 27   d_n = 0+1i 
assign X[4'b0100] [28] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 1^2) * 2^(-2*28) )   n = 28   d_n = 0+1i 
assign X[4'b0100] [29] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 1^2) * 2^(-2*29) )   n = 29   d_n = 0+1i 
assign X[4'b0100] [30] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 1^2) * 2^(-2*30) )   n = 30   d_n = 0+1i 
assign X[4'b0100] [31] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 1^2) * 2^(-2*31) )   n = 31   d_n = 0+1i 
assign X[4'b0100] [32] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 1^2) * 2^(-2*32) )   n = 32   d_n = 0+1i 
assign X[4'b0100] [33] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 1^2) * 2^(-2*33) )   n = 33   d_n = 0+1i 
assign X[4'b0100] [34] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 1^2) * 2^(-2*34) )   n = 34   d_n = 0+1i 
assign X[4'b0100] [35] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 1^2) * 2^(-2*35) )   n = 35   d_n = 0+1i 
assign X[4'b0100] [36] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 1^2) * 2^(-2*36) )   n = 36   d_n = 0+1i 
assign X[4'b0100] [37] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 1^2) * 2^(-2*37) )   n = 37   d_n = 0+1i 
assign X[4'b0100] [38] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 1^2) * 2^(-2*38) )   n = 38   d_n = 0+1i 
assign X[4'b0100] [39] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 1^2) * 2^(-2*39) )   n = 39   d_n = 0+1i 
assign X[4'b0100] [40] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 1^2) * 2^(-2*40) )   n = 40   d_n = 0+1i 
assign X[4'b0100] [41] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 1^2) * 2^(-2*41) )   n = 41   d_n = 0+1i 
assign X[4'b0100] [42] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 1^2) * 2^(-2*42) )   n = 42   d_n = 0+1i 
assign X[4'b0100] [43] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 1^2) * 2^(-2*43) )   n = 43   d_n = 0+1i 
assign X[4'b0100] [44] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 1^2) * 2^(-2*44) )   n = 44   d_n = 0+1i 
assign X[4'b0100] [45] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 1^2) * 2^(-2*45) )   n = 45   d_n = 0+1i 
assign X[4'b0100] [46] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 1^2) * 2^(-2*46) )   n = 46   d_n = 0+1i 
assign X[4'b0100] [47] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 1^2) * 2^(-2*47) )   n = 47   d_n = 0+1i 
assign X[4'b0100] [48] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 1^2) * 2^(-2*48) )   n = 48   d_n = 0+1i 
assign X[4'b0100] [49] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 1^2) * 2^(-2*49) )   n = 49   d_n = 0+1i 
assign X[4'b0100] [50] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 1^2) * 2^(-2*50) )   n = 50   d_n = 0+1i 
assign X[4'b0100] [51] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 1^2) * 2^(-2*51) )   n = 51   d_n = 0+1i 
assign X[4'b0100] [52] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 1^2) * 2^(-2*52) )   n = 52   d_n = 0+1i 
assign X[4'b0100] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 1^2) * 2^(-2*53) )   n = 53   d_n = 0+1i 
assign X[4'b0100] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 1^2) * 2^(-2*54) )   n = 54   d_n = 0+1i 
assign X[4'b0100] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 1^2) * 2^(-2*55) )   n = 55   d_n = 0+1i 
assign X[4'b0100] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 1^2) * 2^(-2*56) )   n = 56   d_n = 0+1i 
assign X[4'b0100] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 1^2) * 2^(-2*57) )   n = 57   d_n = 0+1i 
assign X[4'b0100] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 1^2) * 2^(-2*58) )   n = 58   d_n = 0+1i 
assign X[4'b0100] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 1^2) * 2^(-2*59) )   n = 59   d_n = 0+1i 
assign X[4'b0100] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 1^2) * 2^(-2*60) )   n = 60   d_n = 0+1i 
assign X[4'b0100] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 1^2) * 2^(-2*61) )   n = 61   d_n = 0+1i 
assign X[4'b0100] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 1^2) * 2^(-2*62) )   n = 62   d_n = 0+1i 
assign X[4'b0100] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 1^2) * 2^(-2*63) )   n = 63   d_n = 0+1i 
assign X[4'b0100] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 1^2) * 2^(-2*64) )   n = 64   d_n = 0+1i 
assign X[4'b0101] [01] = 144'h 000000108444104004080420042001020000;  // 0003AA481E1C1C0F20 +0.4581453659370776 = 0.5 * ln( 1 +  1 * 2^(-1+1) + ( 1^2+ 1^2) * 2^(-2*1) )   n =  1   d_n = 1+1i 
assign X[4'b0101] [02] = 144'h 000000040201044100880022020042084400;  // 0001F128F5FAF06EA0 +0.2427539078908503 = 0.5 * ln( 1 +  1 * 2^(-2+1) + ( 1^2+ 1^2) * 2^(-2*2) )   n =  2   d_n = 1+1i 
assign X[4'b0101] [03] = 144'h 000000010008204120108222020402048000;  // 0000FDC8C36AF1F180 +0.1239180819522907 = 0.5 * ln( 1 +  1 * 2^(-3+1) + ( 1^2+ 1^2) * 2^(-2*3) )   n =  3   d_n = 1+1i 
assign X[4'b0101] [04] = 144'h 000000004000220410112040820022220420;  // 00007FB244C76FAB1C +0.0623517392504787 = 0.5 * ln( 1 +  1 * 2^(-4+1) + ( 1^2+ 1^2) * 2^(-2*4) )   n =  4   d_n = 1+1i 
assign X[4'b0101] [05] = 144'h 000000001000008821040412108204480088;  // 00003FF5D2233725F6 +0.0312305848118681 = 0.5 * ln( 1 +  1 * 2^(-5+1) + ( 1^2+ 1^2) * 2^(-2*5) )   n =  5   d_n = 1+1i 
assign X[4'b0101] [06] = 144'h 000000000400000222044101011210441080;  // 00001FFEB291134A38 +0.0156225157283291 = 0.5 * ln( 1 +  1 * 2^(-6+1) + ( 1^2+ 1^2) * 2^(-2*6) )   n =  6   d_n = 1+1i 
assign X[4'b0101] [07] = 144'h 000000000100000008882110404041212102;  // 00000FFFD5D4888CCF +0.0078121858105703 = 0.5 * ln( 1 +  1 * 2^(-7+1) + ( 1^2+ 1^2) * 2^(-2*7) )   n =  7   d_n = 1+1i 
assign X[4'b0101] [08] = 144'h 000000000040000000222204441010101044;  // 000007FFFAB2A4444A +0.0039062104956732 = 0.5 * ln( 1 +  1 * 2^(-8+1) + ( 1^2+ 1^2) * 2^(-2*8) )   n =  8   d_n = 1+1i 
assign X[4'b0101] [09] = 144'h 000000000010000000008888211104040440;  // 000003FFFF55D52228 +0.0019531200474755 = 0.5 * ln( 1 +  1 * 2^(-9+1) + ( 1^2+ 1^2) * 2^(-2*9) )   n =  9   d_n = 1+1i 
assign X[4'b0101] [10] = 144'h 000000000004000000000222220444412101;  // 000001FFFFEAB2A8D1 +0.0009765618800270 = 0.5 * ln( 1 +  1 * 2^(-10+1) + ( 1^2+ 1^2) * 2^(-2*10) )   n = 10   d_n = 1+1i 
assign X[4'b0101] [11] = 144'h 000000000001000000000008888821111044;  // 000000FFFFFD55D54A +0.0004882811724466 = 0.5 * ln( 1 +  1 * 2^(-11+1) + ( 1^2+ 1^2) * 2^(-2*11) )   n = 11   d_n = 1+1i 
assign X[4'b0101] [12] = 144'h 000000000000400000000000222222044444;  // 0000007FFFFFAAB2AA +0.0002441406153023 = 0.5 * ln( 1 +  1 * 2^(-12+1) + ( 1^2+ 1^2) * 2^(-2*12) )   n = 12   d_n = 1+1i 
assign X[4'b0101] [13] = 144'h 000000000000100000000000008888888411;  // 0000003FFFFFF555A5 +0.0001220703112875 = 0.5 * ln( 1 +  1 * 2^(-13+1) + ( 1^2+ 1^2) * 2^(-2*13) )   n = 13   d_n = 1+1i 
assign X[4'b0101] [14] = 144'h 000000000000040000000000000222222200;  // 0000001FFFFFFEAAAF +0.0000610351560984 = 0.5 * ln( 1 +  1 * 2^(-14+1) + ( 1^2+ 1^2) * 2^(-2*14) )   n = 14   d_n = 1+1i 
assign X[4'b0101] [15] = 144'h 000000000000010000000000000008888888;  // 0000000FFFFFFFD555 +0.0000305175781061 = 0.5 * ln( 1 +  1 * 2^(-15+1) + ( 1^2+ 1^2) * 2^(-2*15) )   n = 15   d_n = 1+1i 
assign X[4'b0101] [16] = 144'h 000000000000004000000000000000844444;  // 00000007FFFFFFFAAA +0.0000152587890601 = 0.5 * ln( 1 +  1 * 2^(-16+1) + ( 1^2+ 1^2) * 2^(-2*16) )   n = 16   d_n = 1+1i 
assign X[4'b0101] [17] = 144'h 000000000000001000000000000000021111;  // 00000003FFFFFFFF55 +0.0000076293945310 = 0.5 * ln( 1 +  1 * 2^(-17+1) + ( 1^2+ 1^2) * 2^(-2*17) )   n = 17   d_n = 1+1i 
assign X[4'b0101] [18] = 144'h 000000000000000400000000000000000084;  // 00000001FFFFFFFFFA +0.0000038146972656 = 0.5 * ln( 1 +  1 * 2^(-18+1) + ( 1^2+ 1^2) * 2^(-2*18) )   n = 18   d_n = 1+1i 
assign X[4'b0101] [19] = 144'h 000000000000000100000000000000000002;  // 00000000FFFFFFFFFF +0.0000019073486328 = 0.5 * ln( 1 +  1 * 2^(-19+1) + ( 1^2+ 1^2) * 2^(-2*19) )   n = 19   d_n = 1+1i 
assign X[4'b0101] [20] = 144'h 000000000000000040000000000000000000;  // 000000007FFFFFFFFF +0.0000009536743164 = 0.5 * ln( 1 +  1 * 2^(-20+1) + ( 1^2+ 1^2) * 2^(-2*20) )   n = 20   d_n = 1+1i 
assign X[4'b0101] [21] = 144'h 000000000000000010000000000000000000;  // 000000003FFFFFFFFF +0.0000004768371582 = 0.5 * ln( 1 +  1 * 2^(-21+1) + ( 1^2+ 1^2) * 2^(-2*21) )   n = 21   d_n = 1+1i 
assign X[4'b0101] [22] = 144'h 000000000000000004000000000000000000;  // 000000001FFFFFFFFF +0.0000002384185791 = 0.5 * ln( 1 +  1 * 2^(-22+1) + ( 1^2+ 1^2) * 2^(-2*22) )   n = 22   d_n = 1+1i 
assign X[4'b0101] [23] = 144'h 000000000000000001000000000000000000;  // 000000000FFFFFFFFF +0.0000001192092896 = 0.5 * ln( 1 +  1 * 2^(-23+1) + ( 1^2+ 1^2) * 2^(-2*23) )   n = 23   d_n = 1+1i 
assign X[4'b0101] [24] = 144'h 000000000000000000400000000000000000;  // 0000000007FFFFFFFF +0.0000000596046448 = 0.5 * ln( 1 +  1 * 2^(-24+1) + ( 1^2+ 1^2) * 2^(-2*24) )   n = 24   d_n = 1+1i 
assign X[4'b0101] [25] = 144'h 000000000000000000100000000000000000;  // 0000000003FFFFFFFF +0.0000000298023224 = 0.5 * ln( 1 +  1 * 2^(-25+1) + ( 1^2+ 1^2) * 2^(-2*25) )   n = 25   d_n = 1+1i 
assign X[4'b0101] [26] = 144'h 000000000000000000040000000000002000;  // 0000000001FFFFFFC0 +0.0000000149011611 = 0.5 * ln( 1 +  1 * 2^(-26+1) + ( 1^2+ 1^2) * 2^(-2*26) )   n = 26   d_n = 1+1i 
assign X[4'b0101] [27] = 144'h 000000000000000000010000000000000200;  // 0000000000FFFFFFF0 +0.0000000074505806 = 0.5 * ln( 1 +  1 * 2^(-27+1) + ( 1^2+ 1^2) * 2^(-2*27) )   n = 27   d_n = 1+1i 
assign X[4'b0101] [28] = 144'h 000000000000000000004000000000000020;  // 00000000007FFFFFFC +0.0000000037252903 = 0.5 * ln( 1 +  1 * 2^(-28+1) + ( 1^2+ 1^2) * 2^(-2*28) )   n = 28   d_n = 1+1i 
assign X[4'b0101] [29] = 144'h 000000000000000000001000000000000002;  // 00000000003FFFFFFF +0.0000000018626451 = 0.5 * ln( 1 +  1 * 2^(-29+1) + ( 1^2+ 1^2) * 2^(-2*29) )   n = 29   d_n = 1+1i 
assign X[4'b0101] [30] = 144'h 000000000000000000000400000000000000;  // 00000000001FFFFFFF +0.0000000009313226 = 0.5 * ln( 1 +  1 * 2^(-30+1) + ( 1^2+ 1^2) * 2^(-2*30) )   n = 30   d_n = 1+1i 
assign X[4'b0101] [31] = 144'h 000000000000000000000100000000000000;  // 00000000000FFFFFFF +0.0000000004656613 = 0.5 * ln( 1 +  1 * 2^(-31+1) + ( 1^2+ 1^2) * 2^(-2*31) )   n = 31   d_n = 1+1i 
assign X[4'b0101] [32] = 144'h 000000000000000000000040000000000000;  // 000000000007FFFFFF +0.0000000002328306 = 0.5 * ln( 1 +  1 * 2^(-32+1) + ( 1^2+ 1^2) * 2^(-2*32) )   n = 32   d_n = 1+1i 
assign X[4'b0101] [33] = 144'h 000000000000000000000010000000000000;  // 000000000003FFFFFF +0.0000000001164153 = 0.5 * ln( 1 +  1 * 2^(-33+1) + ( 1^2+ 1^2) * 2^(-2*33) )   n = 33   d_n = 1+1i 
assign X[4'b0101] [34] = 144'h 000000000000000000000004000000000000;  // 000000000001FFFFFF +0.0000000000582077 = 0.5 * ln( 1 +  1 * 2^(-34+1) + ( 1^2+ 1^2) * 2^(-2*34) )   n = 34   d_n = 1+1i 
assign X[4'b0101] [35] = 144'h 000000000000000000000001000000000000;  // 000000000000FFFFFF +0.0000000000291038 = 0.5 * ln( 1 +  1 * 2^(-35+1) + ( 1^2+ 1^2) * 2^(-2*35) )   n = 35   d_n = 1+1i 
assign X[4'b0101] [36] = 144'h 000000000000000000000000400000000000;  // 0000000000007FFFFF +0.0000000000145519 = 0.5 * ln( 1 +  1 * 2^(-36+1) + ( 1^2+ 1^2) * 2^(-2*36) )   n = 36   d_n = 1+1i 
assign X[4'b0101] [37] = 144'h 000000000000000000000000100000000000;  // 0000000000003FFFFF +0.0000000000072760 = 0.5 * ln( 1 +  1 * 2^(-37+1) + ( 1^2+ 1^2) * 2^(-2*37) )   n = 37   d_n = 1+1i 
assign X[4'b0101] [38] = 144'h 000000000000000000000000040000000000;  // 0000000000001FFFFF +0.0000000000036380 = 0.5 * ln( 1 +  1 * 2^(-38+1) + ( 1^2+ 1^2) * 2^(-2*38) )   n = 38   d_n = 1+1i 
assign X[4'b0101] [39] = 144'h 000000000000000000000000010000000000;  // 0000000000000FFFFF +0.0000000000018190 = 0.5 * ln( 1 +  1 * 2^(-39+1) + ( 1^2+ 1^2) * 2^(-2*39) )   n = 39   d_n = 1+1i 
assign X[4'b0101] [40] = 144'h 000000000000000000000000004000000000;  // 00000000000007FFFF +0.0000000000009095 = 0.5 * ln( 1 +  1 * 2^(-40+1) + ( 1^2+ 1^2) * 2^(-2*40) )   n = 40   d_n = 1+1i 
assign X[4'b0101] [41] = 144'h 000000000000000000000000001000000000;  // 00000000000003FFFF +0.0000000000004547 = 0.5 * ln( 1 +  1 * 2^(-41+1) + ( 1^2+ 1^2) * 2^(-2*41) )   n = 41   d_n = 1+1i 
assign X[4'b0101] [42] = 144'h 000000000000000000000000000400000000;  // 00000000000001FFFF +0.0000000000002274 = 0.5 * ln( 1 +  1 * 2^(-42+1) + ( 1^2+ 1^2) * 2^(-2*42) )   n = 42   d_n = 1+1i 
assign X[4'b0101] [43] = 144'h 000000000000000000000000000100000000;  // 00000000000000FFFF +0.0000000000001137 = 0.5 * ln( 1 +  1 * 2^(-43+1) + ( 1^2+ 1^2) * 2^(-2*43) )   n = 43   d_n = 1+1i 
assign X[4'b0101] [44] = 144'h 000000000000000000000000000040000000;  // 000000000000007FFF +0.0000000000000568 = 0.5 * ln( 1 +  1 * 2^(-44+1) + ( 1^2+ 1^2) * 2^(-2*44) )   n = 44   d_n = 1+1i 
assign X[4'b0101] [45] = 144'h 000000000000000000000000000010000000;  // 000000000000003FFF +0.0000000000000284 = 0.5 * ln( 1 +  1 * 2^(-45+1) + ( 1^2+ 1^2) * 2^(-2*45) )   n = 45   d_n = 1+1i 
assign X[4'b0101] [46] = 144'h 000000000000000000000000000004000000;  // 000000000000001FFF +0.0000000000000142 = 0.5 * ln( 1 +  1 * 2^(-46+1) + ( 1^2+ 1^2) * 2^(-2*46) )   n = 46   d_n = 1+1i 
assign X[4'b0101] [47] = 144'h 000000000000000000000000000001000000;  // 000000000000000FFF +0.0000000000000071 = 0.5 * ln( 1 +  1 * 2^(-47+1) + ( 1^2+ 1^2) * 2^(-2*47) )   n = 47   d_n = 1+1i 
assign X[4'b0101] [48] = 144'h 000000000000000000000000000000400000;  // 0000000000000007FF +0.0000000000000036 = 0.5 * ln( 1 +  1 * 2^(-48+1) + ( 1^2+ 1^2) * 2^(-2*48) )   n = 48   d_n = 1+1i 
assign X[4'b0101] [49] = 144'h 000000000000000000000000000000100000;  // 0000000000000003FF +0.0000000000000018 = 0.5 * ln( 1 +  1 * 2^(-49+1) + ( 1^2+ 1^2) * 2^(-2*49) )   n = 49   d_n = 1+1i 
assign X[4'b0101] [50] = 144'h 000000000000000000000000000000040000;  // 0000000000000001FF +0.0000000000000009 = 0.5 * ln( 1 +  1 * 2^(-50+1) + ( 1^2+ 1^2) * 2^(-2*50) )   n = 50   d_n = 1+1i 
assign X[4'b0101] [51] = 144'h 000000000000000000000000000000010000;  // 0000000000000000FF +0.0000000000000004 = 0.5 * ln( 1 +  1 * 2^(-51+1) + ( 1^2+ 1^2) * 2^(-2*51) )   n = 51   d_n = 1+1i 
assign X[4'b0101] [52] = 144'h 000000000000000000000000000000004000;  // 00000000000000007F +0.0000000000000002 = 0.5 * ln( 1 +  1 * 2^(-52+1) + ( 1^2+ 1^2) * 2^(-2*52) )   n = 52   d_n = 1+1i 
assign X[4'b0101] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-53+1) + ( 1^2+ 1^2) * 2^(-2*53) )   n = 53   d_n = 1+1i 
assign X[4'b0101] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-54+1) + ( 1^2+ 1^2) * 2^(-2*54) )   n = 54   d_n = 1+1i 
assign X[4'b0101] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-55+1) + ( 1^2+ 1^2) * 2^(-2*55) )   n = 55   d_n = 1+1i 
assign X[4'b0101] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-56+1) + ( 1^2+ 1^2) * 2^(-2*56) )   n = 56   d_n = 1+1i 
assign X[4'b0101] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-57+1) + ( 1^2+ 1^2) * 2^(-2*57) )   n = 57   d_n = 1+1i 
assign X[4'b0101] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-58+1) + ( 1^2+ 1^2) * 2^(-2*58) )   n = 58   d_n = 1+1i 
assign X[4'b0101] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-59+1) + ( 1^2+ 1^2) * 2^(-2*59) )   n = 59   d_n = 1+1i 
assign X[4'b0101] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-60+1) + ( 1^2+ 1^2) * 2^(-2*60) )   n = 60   d_n = 1+1i 
assign X[4'b0101] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-61+1) + ( 1^2+ 1^2) * 2^(-2*61) )   n = 61   d_n = 1+1i 
assign X[4'b0101] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-62+1) + ( 1^2+ 1^2) * 2^(-2*62) )   n = 62   d_n = 1+1i 
assign X[4'b0101] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-63+1) + ( 1^2+ 1^2) * 2^(-2*63) )   n = 63   d_n = 1+1i 
assign X[4'b0101] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-64+1) + ( 1^2+ 1^2) * 2^(-2*64) )   n = 64   d_n = 1+1i 
assign X[4'b0110] [01] = 144'h 000000010810400020081021211121010400;  // 0000E47FBE3CD4D128 +0.1115717756571049 = 0.5 * ln( 1 +  0 * 2^(-1+1) + ( 0^2+ 1^2) * 2^(-2*1) )   n =  1   d_n = 0+1i 
assign X[4'b0110] [02] = 144'h 000000001008011048048000041220111100;  // 00003E14618022C552 +0.0303123109082174 = 0.5 * ln( 1 +  0 * 2^(-2+1) + ( 0^2+ 1^2) * 2^(-2*2) )   n =  2   d_n = 0+1i 
assign X[4'b0110] [03] = 144'h 000000000100080011104880400800042120;  // 00000FE054587E01CC +0.0077520932679826 = 0.5 * ln( 1 +  0 * 2^(-3+1) + ( 0^2+ 1^2) * 2^(-2*3) )   n =  3   d_n = 0+1i 
assign X[4'b0110] [04] = 144'h 000000000010000800011110488804048404;  // 000003FE01545621A1 +0.0019493202078287 = 0.5 * ln( 1 +  0 * 2^(-4+1) + ( 0^2+ 1^2) * 2^(-2*4) )   n =  4   d_n = 0+1i 
assign X[4'b0110] [05] = 144'h 000000000001000008000011111048888084;  // 000000FFE00554557A +0.0004880429865277 = 0.5 * ln( 1 +  0 * 2^(-5+1) + ( 0^2+ 1^2) * 2^(-2*5) )   n =  5   d_n = 0+1i 
assign X[4'b0110] [06] = 144'h 000000000000100000080000011111100448;  // 0000003FFE00155425 +0.0001220554137636 = 0.5 * ln( 1 +  0 * 2^(-6+1) + ( 0^2+ 1^2) * 2^(-2*6) )   n =  6   d_n = 0+1i 
assign X[4'b0110] [07] = 144'h 000000000000010000000800000011111110;  // 0000000FFFE0005554 +0.0000305166468403 = 0.5 * ln( 1 +  0 * 2^(-7+1) + ( 0^2+ 1^2) * 2^(-2*7) )   n =  7   d_n = 0+1i 
assign X[4'b0110] [08] = 144'h 000000000000001000000008000000011111;  // 00000003FFFE000155 +0.0000076293363242 = 0.5 * ln( 1 +  0 * 2^(-8+1) + ( 0^2+ 1^2) * 2^(-2*8) )   n =  8   d_n = 0+1i 
assign X[4'b0110] [09] = 144'h 000000000000000100000000080000000012;  // 00000000FFFFE00003 +0.0000019073449948 = 0.5 * ln( 1 +  0 * 2^(-9+1) + ( 0^2+ 1^2) * 2^(-2*9) )   n =  9   d_n = 0+1i 
assign X[4'b0110] [10] = 144'h 000000000000000010000000000800000000;  // 000000003FFFFE0000 +0.0000004768369308 = 0.5 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 1^2) * 2^(-2*10) )   n = 10   d_n = 0+1i 
assign X[4'b0110] [11] = 144'h 000000000000000001000000000008000000;  // 000000000FFFFFE000 +0.0000001192092753 = 0.5 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 1^2) * 2^(-2*11) )   n = 11   d_n = 0+1i 
assign X[4'b0110] [12] = 144'h 000000000000000000100000000000080000;  // 0000000003FFFFFE00 +0.0000000298023215 = 0.5 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 1^2) * 2^(-2*12) )   n = 12   d_n = 0+1i 
assign X[4'b0110] [13] = 144'h 000000000000000000010000000000000200;  // 0000000000FFFFFFF0 +0.0000000074505806 = 0.5 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 1^2) * 2^(-2*13) )   n = 13   d_n = 0+1i 
assign X[4'b0110] [14] = 144'h 000000000000000000001000000000000002;  // 00000000003FFFFFFF +0.0000000018626451 = 0.5 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 1^2) * 2^(-2*14) )   n = 14   d_n = 0+1i 
assign X[4'b0110] [15] = 144'h 000000000000000000000100000000000000;  // 00000000000FFFFFFF +0.0000000004656613 = 0.5 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 1^2) * 2^(-2*15) )   n = 15   d_n = 0+1i 
assign X[4'b0110] [16] = 144'h 000000000000000000000010000000000000;  // 000000000003FFFFFF +0.0000000001164153 = 0.5 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 1^2) * 2^(-2*16) )   n = 16   d_n = 0+1i 
assign X[4'b0110] [17] = 144'h 000000000000000000000001000000000000;  // 000000000000FFFFFF +0.0000000000291038 = 0.5 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 1^2) * 2^(-2*17) )   n = 17   d_n = 0+1i 
assign X[4'b0110] [18] = 144'h 000000000000000000000000100000000000;  // 0000000000003FFFFF +0.0000000000072760 = 0.5 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 1^2) * 2^(-2*18) )   n = 18   d_n = 0+1i 
assign X[4'b0110] [19] = 144'h 000000000000000000000000010000000000;  // 0000000000000FFFFF +0.0000000000018190 = 0.5 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 1^2) * 2^(-2*19) )   n = 19   d_n = 0+1i 
assign X[4'b0110] [20] = 144'h 000000000000000000000000001000000000;  // 00000000000003FFFF +0.0000000000004547 = 0.5 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 1^2) * 2^(-2*20) )   n = 20   d_n = 0+1i 
assign X[4'b0110] [21] = 144'h 000000000000000000000000000100000000;  // 00000000000000FFFF +0.0000000000001137 = 0.5 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 1^2) * 2^(-2*21) )   n = 21   d_n = 0+1i 
assign X[4'b0110] [22] = 144'h 000000000000000000000000000010000000;  // 000000000000003FFF +0.0000000000000284 = 0.5 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 1^2) * 2^(-2*22) )   n = 22   d_n = 0+1i 
assign X[4'b0110] [23] = 144'h 000000000000000000000000000001000000;  // 000000000000000FFF +0.0000000000000071 = 0.5 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 1^2) * 2^(-2*23) )   n = 23   d_n = 0+1i 
assign X[4'b0110] [24] = 144'h 000000000000000000000000000000100000;  // 0000000000000003FF +0.0000000000000018 = 0.5 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 1^2) * 2^(-2*24) )   n = 24   d_n = 0+1i 
assign X[4'b0110] [25] = 144'h 000000000000000000000000000000010000;  // 0000000000000000FF +0.0000000000000004 = 0.5 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 1^2) * 2^(-2*25) )   n = 25   d_n = 0+1i 
assign X[4'b0110] [26] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 1^2) * 2^(-2*26) )   n = 26   d_n = 0+1i 
assign X[4'b0110] [27] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 1^2) * 2^(-2*27) )   n = 27   d_n = 0+1i 
assign X[4'b0110] [28] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 1^2) * 2^(-2*28) )   n = 28   d_n = 0+1i 
assign X[4'b0110] [29] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 1^2) * 2^(-2*29) )   n = 29   d_n = 0+1i 
assign X[4'b0110] [30] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 1^2) * 2^(-2*30) )   n = 30   d_n = 0+1i 
assign X[4'b0110] [31] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 1^2) * 2^(-2*31) )   n = 31   d_n = 0+1i 
assign X[4'b0110] [32] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 1^2) * 2^(-2*32) )   n = 32   d_n = 0+1i 
assign X[4'b0110] [33] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 1^2) * 2^(-2*33) )   n = 33   d_n = 0+1i 
assign X[4'b0110] [34] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 1^2) * 2^(-2*34) )   n = 34   d_n = 0+1i 
assign X[4'b0110] [35] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 1^2) * 2^(-2*35) )   n = 35   d_n = 0+1i 
assign X[4'b0110] [36] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 1^2) * 2^(-2*36) )   n = 36   d_n = 0+1i 
assign X[4'b0110] [37] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 1^2) * 2^(-2*37) )   n = 37   d_n = 0+1i 
assign X[4'b0110] [38] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 1^2) * 2^(-2*38) )   n = 38   d_n = 0+1i 
assign X[4'b0110] [39] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 1^2) * 2^(-2*39) )   n = 39   d_n = 0+1i 
assign X[4'b0110] [40] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 1^2) * 2^(-2*40) )   n = 40   d_n = 0+1i 
assign X[4'b0110] [41] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 1^2) * 2^(-2*41) )   n = 41   d_n = 0+1i 
assign X[4'b0110] [42] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 1^2) * 2^(-2*42) )   n = 42   d_n = 0+1i 
assign X[4'b0110] [43] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 1^2) * 2^(-2*43) )   n = 43   d_n = 0+1i 
assign X[4'b0110] [44] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 1^2) * 2^(-2*44) )   n = 44   d_n = 0+1i 
assign X[4'b0110] [45] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 1^2) * 2^(-2*45) )   n = 45   d_n = 0+1i 
assign X[4'b0110] [46] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 1^2) * 2^(-2*46) )   n = 46   d_n = 0+1i 
assign X[4'b0110] [47] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 1^2) * 2^(-2*47) )   n = 47   d_n = 0+1i 
assign X[4'b0110] [48] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 1^2) * 2^(-2*48) )   n = 48   d_n = 0+1i 
assign X[4'b0110] [49] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 1^2) * 2^(-2*49) )   n = 49   d_n = 0+1i 
assign X[4'b0110] [50] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 1^2) * 2^(-2*50) )   n = 50   d_n = 0+1i 
assign X[4'b0110] [51] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 1^2) * 2^(-2*51) )   n = 51   d_n = 0+1i 
assign X[4'b0110] [52] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 1^2) * 2^(-2*52) )   n = 52   d_n = 0+1i 
assign X[4'b0110] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 1^2) * 2^(-2*53) )   n = 53   d_n = 0+1i 
assign X[4'b0110] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 1^2) * 2^(-2*54) )   n = 54   d_n = 0+1i 
assign X[4'b0110] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 1^2) * 2^(-2*55) )   n = 55   d_n = 0+1i 
assign X[4'b0110] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 1^2) * 2^(-2*56) )   n = 56   d_n = 0+1i 
assign X[4'b0110] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 1^2) * 2^(-2*57) )   n = 57   d_n = 0+1i 
assign X[4'b0110] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 1^2) * 2^(-2*58) )   n = 58   d_n = 0+1i 
assign X[4'b0110] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 1^2) * 2^(-2*59) )   n = 59   d_n = 0+1i 
assign X[4'b0110] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 1^2) * 2^(-2*60) )   n = 60   d_n = 0+1i 
assign X[4'b0110] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 1^2) * 2^(-2*61) )   n = 61   d_n = 0+1i 
assign X[4'b0110] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 1^2) * 2^(-2*62) )   n = 62   d_n = 0+1i 
assign X[4'b0110] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 1^2) * 2^(-2*63) )   n = 63   d_n = 0+1i 
assign X[4'b0110] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 1^2) * 2^(-2*64) )   n = 64   d_n = 0+1i 
assign X[4'b0111] [01] = 144'h 000000211084108084000401208120041000;  // FFFD3A37A020B80000 -0.3465735902799726 = 0.5 * ln( 1 + -1 * 2^(-1+1) + (-1^2+ 1^2) * 2^(-2*1) )   n =  1   d_n = -1+1i 
assign X[4'b0111] [02] = 144'h 000000080402208088084808810881121100;  // FFFE1EB75E5D900000 -0.2350018146228677 = 0.5 * ln( 1 + -1 * 2^(-2+1) + (-1^2+ 1^2) * 2^(-2*2) )   n =  2   d_n = -1+1i 
assign X[4'b0111] [03] = 144'h 000000020012108204204484480448101040;  // FFFF03371C9A600000 -0.1234300389657629 = 0.5 * ln( 1 + -1 * 2^(-3+1) + (-1^2+ 1^2) * 2^(-2*3) )   n =  3   d_n = -1+1i 
assign X[4'b0111] [04] = 144'h 000000008000480820220480410044444810;  // FFFF805DBB18900000 -0.0623212226036383 = 0.5 * ln( 1 + -1 * 2^(-4+1) + (-1^2+ 1^2) * 2^(-2*4) )   n =  4   d_n = -1+1i 
assign X[4'b0111] [05] = 144'h 000000002000012212080820444108840110;  // FFFFC00B2DDCA80000 -0.0312286774668733 = 0.5 * ln( 1 + -1 * 2^(-5+1) + (-1^2+ 1^2) * 2^(-2*5) )   n =  5   d_n = -1+1i 
assign X[4'b0111] [06] = 144'h 000000000800000488088202022044888440;  // FFFFE0015D6EF00000 -0.0156223965190538 = 0.5 * ln( 1 + -1 * 2^(-6+1) + (-1^2+ 1^2) * 2^(-2*6) )   n =  6   d_n = -1+1i 
assign X[4'b0111] [07] = 144'h 000000000200000012221220808082120881;  // FFFFF0002B2B780000 -0.0078121783599899 = 0.5 * ln( 1 + -1 * 2^(-7+1) + (-1^2+ 1^2) * 2^(-2*7) )   n =  7   d_n = -1+1i 
assign X[4'b0111] [08] = 144'h 000000000080000000488808882020202088;  // FFFFF800055D580000 -0.0039062100300119 = 0.5 * ln( 1 + -1 * 2^(-8+1) + (-1^2+ 1^2) * 2^(-2*8) )   n =  8   d_n = -1+1i 
assign X[4'b0111] [09] = 144'h 000000000020000000012222122208080810;  // FFFFFC0000AB280000 -0.0019531200183716 = 0.5 * ln( 1 + -1 * 2^(-9+1) + (-1^2+ 1^2) * 2^(-2*9) )   n =  9   d_n = -1+1i 
assign X[4'b0111] [10] = 144'h 000000000008000000000488880888820202;  // FFFFFE000015600000 -0.0009765618782081 = 0.5 * ln( 1 + -1 * 2^(-10+1) + (-1^2+ 1^2) * 2^(-2*10) )   n = 10   d_n = -1+1i 
assign X[4'b0111] [11] = 144'h 000000000002000000000012222212222088;  // FFFFFF000002A80000 -0.0004882811723329 = 0.5 * ln( 1 + -1 * 2^(-11+1) + (-1^2+ 1^2) * 2^(-2*11) )   n = 11   d_n = -1+1i 
assign X[4'b0111] [12] = 144'h 000000000000800000000000488888088888;  // FFFFFF800000580000 -0.0002441406152952 = 0.5 * ln( 1 + -1 * 2^(-12+1) + (-1^2+ 1^2) * 2^(-2*12) )   n = 12   d_n = -1+1i 
assign X[4'b0111] [13] = 144'h 000000000000200000000000012222221022;  // FFFFFFC00000080000 -0.0001220703112871 = 0.5 * ln( 1 + -1 * 2^(-13+1) + (-1^2+ 1^2) * 2^(-2*13) )   n = 13   d_n = -1+1i 
assign X[4'b0111] [14] = 144'h 000000000000080000000000000488888884;  // FFFFFFE00000000000 -0.0000610351560984 = 0.5 * ln( 1 + -1 * 2^(-14+1) + (-1^2+ 1^2) * 2^(-2*14) )   n = 14   d_n = -1+1i 
assign X[4'b0111] [15] = 144'h 000000000000020000000000000012222222;  // FFFFFFF00000000000 -0.0000305175781061 = 0.5 * ln( 1 + -1 * 2^(-15+1) + (-1^2+ 1^2) * 2^(-2*15) )   n = 15   d_n = -1+1i 
assign X[4'b0111] [16] = 144'h 000000000000008000000000000000488888;  // FFFFFFF80000000000 -0.0000152587890601 = 0.5 * ln( 1 + -1 * 2^(-16+1) + (-1^2+ 1^2) * 2^(-2*16) )   n = 16   d_n = -1+1i 
assign X[4'b0111] [17] = 144'h 000000000000002000000000000000012222;  // FFFFFFFC0000000000 -0.0000076293945310 = 0.5 * ln( 1 + -1 * 2^(-17+1) + (-1^2+ 1^2) * 2^(-2*17) )   n = 17   d_n = -1+1i 
assign X[4'b0111] [18] = 144'h 000000000000000800000000000000000048;  // FFFFFFFE0000000000 -0.0000038146972656 = 0.5 * ln( 1 + -1 * 2^(-18+1) + (-1^2+ 1^2) * 2^(-2*18) )   n = 18   d_n = -1+1i 
assign X[4'b0111] [19] = 144'h 000000000000000200000000000000000001;  // FFFFFFFF0000000000 -0.0000019073486328 = 0.5 * ln( 1 + -1 * 2^(-19+1) + (-1^2+ 1^2) * 2^(-2*19) )   n = 19   d_n = -1+1i 
assign X[4'b0111] [20] = 144'h 000000000000000080000000000000000000;  // FFFFFFFF8000000000 -0.0000009536743164 = 0.5 * ln( 1 + -1 * 2^(-20+1) + (-1^2+ 1^2) * 2^(-2*20) )   n = 20   d_n = -1+1i 
assign X[4'b0111] [21] = 144'h 000000000000000020000000000000000000;  // FFFFFFFFC000000000 -0.0000004768371582 = 0.5 * ln( 1 + -1 * 2^(-21+1) + (-1^2+ 1^2) * 2^(-2*21) )   n = 21   d_n = -1+1i 
assign X[4'b0111] [22] = 144'h 000000000000000008000000000000000000;  // FFFFFFFFE000000000 -0.0000002384185791 = 0.5 * ln( 1 + -1 * 2^(-22+1) + (-1^2+ 1^2) * 2^(-2*22) )   n = 22   d_n = -1+1i 
assign X[4'b0111] [23] = 144'h 000000000000000002000000000000000000;  // FFFFFFFFF000000000 -0.0000001192092896 = 0.5 * ln( 1 + -1 * 2^(-23+1) + (-1^2+ 1^2) * 2^(-2*23) )   n = 23   d_n = -1+1i 
assign X[4'b0111] [24] = 144'h 000000000000000000800000000000000000;  // FFFFFFFFF800000000 -0.0000000596046448 = 0.5 * ln( 1 + -1 * 2^(-24+1) + (-1^2+ 1^2) * 2^(-2*24) )   n = 24   d_n = -1+1i 
assign X[4'b0111] [25] = 144'h 000000000000000000200000000000000000;  // FFFFFFFFFC00000000 -0.0000000298023224 = 0.5 * ln( 1 + -1 * 2^(-25+1) + (-1^2+ 1^2) * 2^(-2*25) )   n = 25   d_n = -1+1i 
assign X[4'b0111] [26] = 144'h 000000000000000000080000000000000000;  // FFFFFFFFFE00000000 -0.0000000149011612 = 0.5 * ln( 1 + -1 * 2^(-26+1) + (-1^2+ 1^2) * 2^(-2*26) )   n = 26   d_n = -1+1i 
assign X[4'b0111] [27] = 144'h 000000000000000000020000000000000200;  // FFFFFFFFFF00000000 -0.0000000074505806 = 0.5 * ln( 1 + -1 * 2^(-27+1) + (-1^2+ 1^2) * 2^(-2*27) )   n = 27   d_n = -1+1i 
assign X[4'b0111] [28] = 144'h 000000000000000000008000000000000020;  // FFFFFFFFFF80000000 -0.0000000037252903 = 0.5 * ln( 1 + -1 * 2^(-28+1) + (-1^2+ 1^2) * 2^(-2*28) )   n = 28   d_n = -1+1i 
assign X[4'b0111] [29] = 144'h 000000000000000000002000000000000002;  // FFFFFFFFFFC0000000 -0.0000000018626452 = 0.5 * ln( 1 + -1 * 2^(-29+1) + (-1^2+ 1^2) * 2^(-2*29) )   n = 29   d_n = -1+1i 
assign X[4'b0111] [30] = 144'h 000000000000000000000800000000000000;  // FFFFFFFFFFE0000000 -0.0000000009313226 = 0.5 * ln( 1 + -1 * 2^(-30+1) + (-1^2+ 1^2) * 2^(-2*30) )   n = 30   d_n = -1+1i 
assign X[4'b0111] [31] = 144'h 000000000000000000000200000000000000;  // FFFFFFFFFFF0000000 -0.0000000004656613 = 0.5 * ln( 1 + -1 * 2^(-31+1) + (-1^2+ 1^2) * 2^(-2*31) )   n = 31   d_n = -1+1i 
assign X[4'b0111] [32] = 144'h 000000000000000000000080000000000000;  // FFFFFFFFFFF8000000 -0.0000000002328306 = 0.5 * ln( 1 + -1 * 2^(-32+1) + (-1^2+ 1^2) * 2^(-2*32) )   n = 32   d_n = -1+1i 
assign X[4'b0111] [33] = 144'h 000000000000000000000020000000000000;  // FFFFFFFFFFFC000000 -0.0000000001164153 = 0.5 * ln( 1 + -1 * 2^(-33+1) + (-1^2+ 1^2) * 2^(-2*33) )   n = 33   d_n = -1+1i 
assign X[4'b0111] [34] = 144'h 000000000000000000000008000000000000;  // FFFFFFFFFFFE000000 -0.0000000000582077 = 0.5 * ln( 1 + -1 * 2^(-34+1) + (-1^2+ 1^2) * 2^(-2*34) )   n = 34   d_n = -1+1i 
assign X[4'b0111] [35] = 144'h 000000000000000000000002000000000000;  // FFFFFFFFFFFF000000 -0.0000000000291038 = 0.5 * ln( 1 + -1 * 2^(-35+1) + (-1^2+ 1^2) * 2^(-2*35) )   n = 35   d_n = -1+1i 
assign X[4'b0111] [36] = 144'h 000000000000000000000000800000000000;  // FFFFFFFFFFFF800000 -0.0000000000145519 = 0.5 * ln( 1 + -1 * 2^(-36+1) + (-1^2+ 1^2) * 2^(-2*36) )   n = 36   d_n = -1+1i 
assign X[4'b0111] [37] = 144'h 000000000000000000000000200000000000;  // FFFFFFFFFFFFC00000 -0.0000000000072760 = 0.5 * ln( 1 + -1 * 2^(-37+1) + (-1^2+ 1^2) * 2^(-2*37) )   n = 37   d_n = -1+1i 
assign X[4'b0111] [38] = 144'h 000000000000000000000000080000000000;  // FFFFFFFFFFFFE00000 -0.0000000000036380 = 0.5 * ln( 1 + -1 * 2^(-38+1) + (-1^2+ 1^2) * 2^(-2*38) )   n = 38   d_n = -1+1i 
assign X[4'b0111] [39] = 144'h 000000000000000000000000020000000000;  // FFFFFFFFFFFFF00000 -0.0000000000018190 = 0.5 * ln( 1 + -1 * 2^(-39+1) + (-1^2+ 1^2) * 2^(-2*39) )   n = 39   d_n = -1+1i 
assign X[4'b0111] [40] = 144'h 000000000000000000000000008000000000;  // FFFFFFFFFFFFF80000 -0.0000000000009095 = 0.5 * ln( 1 + -1 * 2^(-40+1) + (-1^2+ 1^2) * 2^(-2*40) )   n = 40   d_n = -1+1i 
assign X[4'b0111] [41] = 144'h 000000000000000000000000002000000000;  // FFFFFFFFFFFFF80000 -0.0000000000004547 = 0.5 * ln( 1 + -1 * 2^(-41+1) + (-1^2+ 1^2) * 2^(-2*41) )   n = 41   d_n = -1+1i 
assign X[4'b0111] [42] = 144'h 000000000000000000000000000800000000;  // 1000000000000000000 -0.0000000000002274 = 0.5 * ln( 1 + -1 * 2^(-42+1) + (-1^2+ 1^2) * 2^(-2*42) )   n = 42   d_n = -1+1i 
assign X[4'b0111] [43] = 144'h 000000000000000000000000000200000000;  // 1000000000000000000 -0.0000000000001137 = 0.5 * ln( 1 + -1 * 2^(-43+1) + (-1^2+ 1^2) * 2^(-2*43) )   n = 43   d_n = -1+1i 
assign X[4'b0111] [44] = 144'h 000000000000000000000000000080000000;  // 1000000000000000000 -0.0000000000000568 = 0.5 * ln( 1 + -1 * 2^(-44+1) + (-1^2+ 1^2) * 2^(-2*44) )   n = 44   d_n = -1+1i 
assign X[4'b0111] [45] = 144'h 000000000000000000000000000020000000;  // 1000000000000000000 -0.0000000000000284 = 0.5 * ln( 1 + -1 * 2^(-45+1) + (-1^2+ 1^2) * 2^(-2*45) )   n = 45   d_n = -1+1i 
assign X[4'b0111] [46] = 144'h 000000000000000000000000000008000000;  // 1000000000000000000 -0.0000000000000142 = 0.5 * ln( 1 + -1 * 2^(-46+1) + (-1^2+ 1^2) * 2^(-2*46) )   n = 46   d_n = -1+1i 
assign X[4'b0111] [47] = 144'h 000000000000000000000000000002000000;  // 1000000000000000000 -0.0000000000000071 = 0.5 * ln( 1 + -1 * 2^(-47+1) + (-1^2+ 1^2) * 2^(-2*47) )   n = 47   d_n = -1+1i 
assign X[4'b0111] [48] = 144'h 000000000000000000000000000000800000;  // 1000000000000000000 -0.0000000000000036 = 0.5 * ln( 1 + -1 * 2^(-48+1) + (-1^2+ 1^2) * 2^(-2*48) )   n = 48   d_n = -1+1i 
assign X[4'b0111] [49] = 144'h 000000000000000000000000000000200000;  // 1000000000000000000 -0.0000000000000018 = 0.5 * ln( 1 + -1 * 2^(-49+1) + (-1^2+ 1^2) * 2^(-2*49) )   n = 49   d_n = -1+1i 
assign X[4'b0111] [50] = 144'h 000000000000000000000000000000080000;  // 1000000000000000000 -0.0000000000000009 = 0.5 * ln( 1 + -1 * 2^(-50+1) + (-1^2+ 1^2) * 2^(-2*50) )   n = 50   d_n = -1+1i 
assign X[4'b0111] [51] = 144'h 000000000000000000000000000000020000;  // 1000000000000000000 -0.0000000000000004 = 0.5 * ln( 1 + -1 * 2^(-51+1) + (-1^2+ 1^2) * 2^(-2*51) )   n = 51   d_n = -1+1i 
assign X[4'b0111] [52] = 144'h 000000000000000000000000000000008000;  // 1000000000000000000 -0.0000000000000002 = 0.5 * ln( 1 + -1 * 2^(-52+1) + (-1^2+ 1^2) * 2^(-2*52) )   n = 52   d_n = -1+1i 
assign X[4'b0111] [53] = 144'h 000000000000000000000000000000002000;  // 1000000000000000000 -0.0000000000000001 = 0.5 * ln( 1 + -1 * 2^(-53+1) + (-1^2+ 1^2) * 2^(-2*53) )   n = 53   d_n = -1+1i 
assign X[4'b0111] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-54+1) + (-1^2+ 1^2) * 2^(-2*54) )   n = 54   d_n = -1+1i 
assign X[4'b0111] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-55+1) + (-1^2+ 1^2) * 2^(-2*55) )   n = 55   d_n = -1+1i 
assign X[4'b0111] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-56+1) + (-1^2+ 1^2) * 2^(-2*56) )   n = 56   d_n = -1+1i 
assign X[4'b0111] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-57+1) + (-1^2+ 1^2) * 2^(-2*57) )   n = 57   d_n = -1+1i 
assign X[4'b0111] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-58+1) + (-1^2+ 1^2) * 2^(-2*58) )   n = 58   d_n = -1+1i 
assign X[4'b0111] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-59+1) + (-1^2+ 1^2) * 2^(-2*59) )   n = 59   d_n = -1+1i 
assign X[4'b0111] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-60+1) + (-1^2+ 1^2) * 2^(-2*60) )   n = 60   d_n = -1+1i 
assign X[4'b0111] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-61+1) + (-1^2+ 1^2) * 2^(-2*61) )   n = 61   d_n = -1+1i 
assign X[4'b0111] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-62+1) + (-1^2+ 1^2) * 2^(-2*62) )   n = 62   d_n = -1+1i 
assign X[4'b0111] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-63+1) + (-1^2+ 1^2) * 2^(-2*63) )   n = 63   d_n = -1+1i 
assign X[4'b0111] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-64+1) + (-1^2+ 1^2) * 2^(-2*64) )   n = 64   d_n = -1+1i 
assign X[4'b1000] [01] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-1+1) + ( 0^2+ 0^2) * 2^(-2*1) )   n =  1   d_n = 0 
assign X[4'b1000] [02] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-2+1) + ( 0^2+ 0^2) * 2^(-2*2) )   n =  2   d_n = 0 
assign X[4'b1000] [03] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-3+1) + ( 0^2+ 0^2) * 2^(-2*3) )   n =  3   d_n = 0 
assign X[4'b1000] [04] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-4+1) + ( 0^2+ 0^2) * 2^(-2*4) )   n =  4   d_n = 0 
assign X[4'b1000] [05] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-5+1) + ( 0^2+ 0^2) * 2^(-2*5) )   n =  5   d_n = 0 
assign X[4'b1000] [06] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-6+1) + ( 0^2+ 0^2) * 2^(-2*6) )   n =  6   d_n = 0 
assign X[4'b1000] [07] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-7+1) + ( 0^2+ 0^2) * 2^(-2*7) )   n =  7   d_n = 0 
assign X[4'b1000] [08] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-8+1) + ( 0^2+ 0^2) * 2^(-2*8) )   n =  8   d_n = 0 
assign X[4'b1000] [09] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-9+1) + ( 0^2+ 0^2) * 2^(-2*9) )   n =  9   d_n = 0 
assign X[4'b1000] [10] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = 0 
assign X[4'b1000] [11] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = 0 
assign X[4'b1000] [12] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = 0 
assign X[4'b1000] [13] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = 0 
assign X[4'b1000] [14] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = 0 
assign X[4'b1000] [15] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = 0 
assign X[4'b1000] [16] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = 0 
assign X[4'b1000] [17] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = 0 
assign X[4'b1000] [18] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = 0 
assign X[4'b1000] [19] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = 0 
assign X[4'b1000] [20] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = 0 
assign X[4'b1000] [21] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = 0 
assign X[4'b1000] [22] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = 0 
assign X[4'b1000] [23] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = 0 
assign X[4'b1000] [24] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = 0 
assign X[4'b1000] [25] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = 0 
assign X[4'b1000] [26] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = 0 
assign X[4'b1000] [27] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = 0 
assign X[4'b1000] [28] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = 0 
assign X[4'b1000] [29] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = 0 
assign X[4'b1000] [30] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = 0 
assign X[4'b1000] [31] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = 0 
assign X[4'b1000] [32] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = 0 
assign X[4'b1000] [33] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = 0 
assign X[4'b1000] [34] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = 0 
assign X[4'b1000] [35] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = 0 
assign X[4'b1000] [36] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = 0 
assign X[4'b1000] [37] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = 0 
assign X[4'b1000] [38] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = 0 
assign X[4'b1000] [39] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = 0 
assign X[4'b1000] [40] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = 0 
assign X[4'b1000] [41] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = 0 
assign X[4'b1000] [42] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = 0 
assign X[4'b1000] [43] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = 0 
assign X[4'b1000] [44] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = 0 
assign X[4'b1000] [45] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = 0 
assign X[4'b1000] [46] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = 0 
assign X[4'b1000] [47] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = 0 
assign X[4'b1000] [48] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = 0 
assign X[4'b1000] [49] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = 0 
assign X[4'b1000] [50] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = 0 
assign X[4'b1000] [51] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = 0 
assign X[4'b1000] [52] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = 0 
assign X[4'b1000] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = 0 
assign X[4'b1000] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = 0 
assign X[4'b1000] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = 0 
assign X[4'b1000] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = 0 
assign X[4'b1000] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = 0 
assign X[4'b1000] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = 0 
assign X[4'b1000] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = 0 
assign X[4'b1000] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = 0 
assign X[4'b1000] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = 0 
assign X[4'b1000] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = 0 
assign X[4'b1000] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = 0 
assign X[4'b1000] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = 0 
assign X[4'b1001] [01] = 144'h 000000121008481040088480021200448000;  // 00033E647D97F30980 +0.4054651081081644 = 0.5 * ln( 1 +  1 * 2^(-1+1) + ( 1^2+ 0^2) * 2^(-2*1) )   n =  1   d_n = 1 
assign X[4'b1001] [02] = 144'h 000000042041000080204084844484040400;  // 0001C8FF7C79A9A220 +0.2231435513142098 = 0.5 * ln( 1 +  1 * 2^(-2+1) + ( 1^2+ 0^2) * 2^(-2*2) )   n =  2   d_n = 1 
assign X[4'b1001] [03] = 144'h 000000010201108010208204888084821200;  // 0000F1383B71579730 +0.1177830356563835 = 0.5 * ln( 1 +  1 * 2^(-3+1) + ( 1^2+ 0^2) * 2^(-2*3) )   n =  3   d_n = 1 
assign X[4'b1001] [04] = 144'h 000000004020044120120000104880444480;  // 00007C28C300458A98 +0.0606246218164348 = 0.5 * ln( 1 +  1 * 2^(-4+1) + ( 1^2+ 0^2) * 2^(-2*4) )   n =  4   d_n = 1 
assign X[4'b1001] [05] = 144'h 000000001002001110880421020048480000;  // 00003F05361CF06600 +0.0307716586667537 = 0.5 * ln( 1 +  1 * 2^(-5+1) + ( 1^2+ 0^2) * 2^(-2*5) )   n =  5   d_n = 1 
assign X[4'b1001] [06] = 144'h 000000000400200044412201002000100810;  // 00001FC0A8B0FC03E4 +0.0155041865359653 = 0.5 * ln( 1 +  1 * 2^(-6+1) + ( 1^2+ 0^2) * 2^(-2*6) )   n =  6   d_n = 1 
assign X[4'b1001] [07] = 144'h 000000000100020001111088804012102010;  // 00000FF015358833C4 +0.0077821404420549 = 0.5 * ln( 1 +  1 * 2^(-7+1) + ( 1^2+ 0^2) * 2^(-2*7) )   n =  7   d_n = 1 
assign X[4'b1001] [08] = 144'h 000000000040002000044441222010120200;  // 000007FC02A8AC42F0 +0.0038986404156573 = 0.5 * ln( 1 +  1 * 2^(-8+1) + ( 1^2+ 0^2) * 2^(-2*8) )   n =  8   d_n = 1 
assign X[4'b1001] [09] = 144'h 000000000010000200001111108888040421;  // 000003FF005535621C +0.0019512201312617 = 0.5 * ln( 1 +  1 * 2^(-9+1) + ( 1^2+ 0^2) * 2^(-2*9) )   n =  9   d_n = 1 
assign X[4'b1001] [10] = 144'h 000000000004000020000044444122220101;  // 000001FFC00AA8AB11 +0.0009760859730555 = 0.5 * ln( 1 +  1 * 2^(-10+1) + ( 1^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = 1 
assign X[4'b1001] [11] = 144'h 000000000001000002000001111110888880;  // 000000FFF001553558 +0.0004881620795014 = 0.5 * ln( 1 +  1 * 2^(-11+1) + ( 1^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = 1 
assign X[4'b1001] [12] = 144'h 000000000000400000200000044444412222;  // 0000007FFC002AA8AA +0.0002441108275274 = 0.5 * ln( 1 +  1 * 2^(-12+1) + ( 1^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = 1 
assign X[4'b1001] [13] = 144'h 000000000000100000020000001111111211;  // 0000003FFF00055535 +0.0001220628625257 = 0.5 * ln( 1 +  1 * 2^(-13+1) + ( 1^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = 1 
assign X[4'b1001] [14] = 144'h 000000000000040000002000000044444440;  // 0000001FFFC000AAA8 +0.0000610332936806 = 0.5 * ln( 1 +  1 * 2^(-14+1) + ( 1^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = 1 
assign X[4'b1001] [15] = 144'h 000000000000010000000200000001111111;  // 0000000FFFF0001555 +0.0000305171124732 = 0.5 * ln( 1 +  1 * 2^(-15+1) + ( 1^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = 1 
assign X[4'b1001] [16] = 144'h 000000000000004000000020000000044444;  // 00000007FFFC0002AA +0.0000152586726484 = 0.5 * ln( 1 +  1 * 2^(-16+1) + ( 1^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = 1 
assign X[4'b1001] [17] = 144'h 000000000000001000000002000000001111;  // 00000003FFFF000055 +0.0000076293654276 = 0.5 * ln( 1 +  1 * 2^(-17+1) + ( 1^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = 1 
assign X[4'b1001] [18] = 144'h 000000000000000400000000200000000044;  // 00000001FFFFC0000A +0.0000038146899897 = 0.5 * ln( 1 +  1 * 2^(-18+1) + ( 1^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = 1 
assign X[4'b1001] [19] = 144'h 000000000000000100000000020000000001;  // 00000000FFFFF00001 +0.0000019073468138 = 0.5 * ln( 1 +  1 * 2^(-19+1) + ( 1^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = 1 
assign X[4'b1001] [20] = 144'h 000000000000000040000000002000000000;  // 000000007FFFFC0000 +0.0000009536738617 = 0.5 * ln( 1 +  1 * 2^(-20+1) + ( 1^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = 1 
assign X[4'b1001] [21] = 144'h 000000000000000010000000000200000000;  // 000000003FFFFF0000 +0.0000004768370445 = 0.5 * ln( 1 +  1 * 2^(-21+1) + ( 1^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = 1 
assign X[4'b1001] [22] = 144'h 000000000000000004000000000020000000;  // 000000001FFFFFC000 +0.0000002384185507 = 0.5 * ln( 1 +  1 * 2^(-22+1) + ( 1^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = 1 
assign X[4'b1001] [23] = 144'h 000000000000000001000000000002000000;  // 000000000FFFFFF000 +0.0000001192092824 = 0.5 * ln( 1 +  1 * 2^(-23+1) + ( 1^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = 1 
assign X[4'b1001] [24] = 144'h 000000000000000000400000000000200000;  // 0000000007FFFFFC00 +0.0000000596046430 = 0.5 * ln( 1 +  1 * 2^(-24+1) + ( 1^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = 1 
assign X[4'b1001] [25] = 144'h 000000000000000000100000000000020000;  // 0000000003FFFFFF00 +0.0000000298023219 = 0.5 * ln( 1 +  1 * 2^(-25+1) + ( 1^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = 1 
assign X[4'b1001] [26] = 144'h 000000000000000000040000000000002000;  // 0000000001FFFFFFC0 +0.0000000149011611 = 0.5 * ln( 1 +  1 * 2^(-26+1) + ( 1^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = 1 
assign X[4'b1001] [27] = 144'h 000000000000000000010000000000000200;  // 0000000000FFFFFFF0 +0.0000000074505806 = 0.5 * ln( 1 +  1 * 2^(-27+1) + ( 1^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = 1 
assign X[4'b1001] [28] = 144'h 000000000000000000004000000000000020;  // 00000000007FFFFFFC +0.0000000037252903 = 0.5 * ln( 1 +  1 * 2^(-28+1) + ( 1^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = 1 
assign X[4'b1001] [29] = 144'h 000000000000000000001000000000000002;  // 00000000003FFFFFFF +0.0000000018626451 = 0.5 * ln( 1 +  1 * 2^(-29+1) + ( 1^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = 1 
assign X[4'b1001] [30] = 144'h 000000000000000000000400000000000000;  // 00000000001FFFFFFF +0.0000000009313226 = 0.5 * ln( 1 +  1 * 2^(-30+1) + ( 1^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = 1 
assign X[4'b1001] [31] = 144'h 000000000000000000000100000000000000;  // 00000000000FFFFFFF +0.0000000004656613 = 0.5 * ln( 1 +  1 * 2^(-31+1) + ( 1^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = 1 
assign X[4'b1001] [32] = 144'h 000000000000000000000040000000000000;  // 000000000007FFFFFF +0.0000000002328306 = 0.5 * ln( 1 +  1 * 2^(-32+1) + ( 1^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = 1 
assign X[4'b1001] [33] = 144'h 000000000000000000000010000000000000;  // 000000000003FFFFFF +0.0000000001164153 = 0.5 * ln( 1 +  1 * 2^(-33+1) + ( 1^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = 1 
assign X[4'b1001] [34] = 144'h 000000000000000000000004000000000000;  // 000000000001FFFFFF +0.0000000000582077 = 0.5 * ln( 1 +  1 * 2^(-34+1) + ( 1^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = 1 
assign X[4'b1001] [35] = 144'h 000000000000000000000001000000000000;  // 000000000000FFFFFF +0.0000000000291038 = 0.5 * ln( 1 +  1 * 2^(-35+1) + ( 1^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = 1 
assign X[4'b1001] [36] = 144'h 000000000000000000000000400000000000;  // 0000000000007FFFFF +0.0000000000145519 = 0.5 * ln( 1 +  1 * 2^(-36+1) + ( 1^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = 1 
assign X[4'b1001] [37] = 144'h 000000000000000000000000100000000000;  // 0000000000003FFFFF +0.0000000000072760 = 0.5 * ln( 1 +  1 * 2^(-37+1) + ( 1^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = 1 
assign X[4'b1001] [38] = 144'h 000000000000000000000000040000000000;  // 0000000000001FFFFF +0.0000000000036380 = 0.5 * ln( 1 +  1 * 2^(-38+1) + ( 1^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = 1 
assign X[4'b1001] [39] = 144'h 000000000000000000000000010000000000;  // 0000000000000FFFFF +0.0000000000018190 = 0.5 * ln( 1 +  1 * 2^(-39+1) + ( 1^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = 1 
assign X[4'b1001] [40] = 144'h 000000000000000000000000004000000000;  // 00000000000007FFFF +0.0000000000009095 = 0.5 * ln( 1 +  1 * 2^(-40+1) + ( 1^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = 1 
assign X[4'b1001] [41] = 144'h 000000000000000000000000001000000000;  // 00000000000003FFFF +0.0000000000004547 = 0.5 * ln( 1 +  1 * 2^(-41+1) + ( 1^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = 1 
assign X[4'b1001] [42] = 144'h 000000000000000000000000000400000000;  // 00000000000001FFFF +0.0000000000002274 = 0.5 * ln( 1 +  1 * 2^(-42+1) + ( 1^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = 1 
assign X[4'b1001] [43] = 144'h 000000000000000000000000000100000000;  // 00000000000000FFFF +0.0000000000001137 = 0.5 * ln( 1 +  1 * 2^(-43+1) + ( 1^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = 1 
assign X[4'b1001] [44] = 144'h 000000000000000000000000000040000000;  // 000000000000007FFF +0.0000000000000568 = 0.5 * ln( 1 +  1 * 2^(-44+1) + ( 1^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = 1 
assign X[4'b1001] [45] = 144'h 000000000000000000000000000010000000;  // 000000000000003FFF +0.0000000000000284 = 0.5 * ln( 1 +  1 * 2^(-45+1) + ( 1^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = 1 
assign X[4'b1001] [46] = 144'h 000000000000000000000000000004000000;  // 000000000000001FFF +0.0000000000000142 = 0.5 * ln( 1 +  1 * 2^(-46+1) + ( 1^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = 1 
assign X[4'b1001] [47] = 144'h 000000000000000000000000000001000000;  // 000000000000000FFF +0.0000000000000071 = 0.5 * ln( 1 +  1 * 2^(-47+1) + ( 1^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = 1 
assign X[4'b1001] [48] = 144'h 000000000000000000000000000000400000;  // 0000000000000007FF +0.0000000000000036 = 0.5 * ln( 1 +  1 * 2^(-48+1) + ( 1^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = 1 
assign X[4'b1001] [49] = 144'h 000000000000000000000000000000100000;  // 0000000000000003FF +0.0000000000000018 = 0.5 * ln( 1 +  1 * 2^(-49+1) + ( 1^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = 1 
assign X[4'b1001] [50] = 144'h 000000000000000000000000000000040000;  // 0000000000000001FF +0.0000000000000009 = 0.5 * ln( 1 +  1 * 2^(-50+1) + ( 1^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = 1 
assign X[4'b1001] [51] = 144'h 000000000000000000000000000000010000;  // 0000000000000000FF +0.0000000000000004 = 0.5 * ln( 1 +  1 * 2^(-51+1) + ( 1^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = 1 
assign X[4'b1001] [52] = 144'h 000000000000000000000000000000004000;  // 00000000000000007F +0.0000000000000002 = 0.5 * ln( 1 +  1 * 2^(-52+1) + ( 1^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = 1 
assign X[4'b1001] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-53+1) + ( 1^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = 1 
assign X[4'b1001] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-54+1) + ( 1^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = 1 
assign X[4'b1001] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-55+1) + ( 1^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = 1 
assign X[4'b1001] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-56+1) + ( 1^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = 1 
assign X[4'b1001] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-57+1) + ( 1^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = 1 
assign X[4'b1001] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-58+1) + ( 1^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = 1 
assign X[4'b1001] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-59+1) + ( 1^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = 1 
assign X[4'b1001] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-60+1) + ( 1^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = 1 
assign X[4'b1001] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-61+1) + ( 1^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = 1 
assign X[4'b1001] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-62+1) + ( 1^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = 1 
assign X[4'b1001] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-63+1) + ( 1^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = 1 
assign X[4'b1001] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-64+1) + ( 1^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = 1 
assign X[4'b1010] [01] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-1+1) + ( 0^2+ 0^2) * 2^(-2*1) )   n =  1   d_n = -0 
assign X[4'b1010] [02] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-2+1) + ( 0^2+ 0^2) * 2^(-2*2) )   n =  2   d_n = -0 
assign X[4'b1010] [03] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-3+1) + ( 0^2+ 0^2) * 2^(-2*3) )   n =  3   d_n = -0 
assign X[4'b1010] [04] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-4+1) + ( 0^2+ 0^2) * 2^(-2*4) )   n =  4   d_n = -0 
assign X[4'b1010] [05] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-5+1) + ( 0^2+ 0^2) * 2^(-2*5) )   n =  5   d_n = -0 
assign X[4'b1010] [06] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-6+1) + ( 0^2+ 0^2) * 2^(-2*6) )   n =  6   d_n = -0 
assign X[4'b1010] [07] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-7+1) + ( 0^2+ 0^2) * 2^(-2*7) )   n =  7   d_n = -0 
assign X[4'b1010] [08] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-8+1) + ( 0^2+ 0^2) * 2^(-2*8) )   n =  8   d_n = -0 
assign X[4'b1010] [09] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-9+1) + ( 0^2+ 0^2) * 2^(-2*9) )   n =  9   d_n = -0 
assign X[4'b1010] [10] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = -0 
assign X[4'b1010] [11] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = -0 
assign X[4'b1010] [12] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = -0 
assign X[4'b1010] [13] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = -0 
assign X[4'b1010] [14] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = -0 
assign X[4'b1010] [15] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = -0 
assign X[4'b1010] [16] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = -0 
assign X[4'b1010] [17] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = -0 
assign X[4'b1010] [18] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = -0 
assign X[4'b1010] [19] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = -0 
assign X[4'b1010] [20] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = -0 
assign X[4'b1010] [21] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = -0 
assign X[4'b1010] [22] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = -0 
assign X[4'b1010] [23] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = -0 
assign X[4'b1010] [24] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = -0 
assign X[4'b1010] [25] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = -0 
assign X[4'b1010] [26] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = -0 
assign X[4'b1010] [27] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = -0 
assign X[4'b1010] [28] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = -0 
assign X[4'b1010] [29] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = -0 
assign X[4'b1010] [30] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = -0 
assign X[4'b1010] [31] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = -0 
assign X[4'b1010] [32] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = -0 
assign X[4'b1010] [33] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = -0 
assign X[4'b1010] [34] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = -0 
assign X[4'b1010] [35] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = -0 
assign X[4'b1010] [36] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = -0 
assign X[4'b1010] [37] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = -0 
assign X[4'b1010] [38] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = -0 
assign X[4'b1010] [39] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = -0 
assign X[4'b1010] [40] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = -0 
assign X[4'b1010] [41] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = -0 
assign X[4'b1010] [42] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = -0 
assign X[4'b1010] [43] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = -0 
assign X[4'b1010] [44] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = -0 
assign X[4'b1010] [45] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = -0 
assign X[4'b1010] [46] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = -0 
assign X[4'b1010] [47] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = -0 
assign X[4'b1010] [48] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = -0 
assign X[4'b1010] [49] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = -0 
assign X[4'b1010] [50] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = -0 
assign X[4'b1010] [51] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = -0 
assign X[4'b1010] [52] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = -0 
assign X[4'b1010] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = -0 
assign X[4'b1010] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = -0 
assign X[4'b1010] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = -0 
assign X[4'b1010] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = -0 
assign X[4'b1010] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = -0 
assign X[4'b1010] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = -0 
assign X[4'b1010] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = -0 
assign X[4'b1010] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = -0 
assign X[4'b1010] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = -0 
assign X[4'b1010] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = -0 
assign X[4'b1010] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = -0 
assign X[4'b1010] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = -0 
assign X[4'b1011] [01] = 144'h 000000844210420210001004820480101000;  // FFFA746F4041700000 -0.6931471805599453 = 0.5 * ln( 1 + -1 * 2^(-1+1) + (-1^2+ 0^2) * 2^(-2*1) )   n =  1   d_n = -1 
assign X[4'b1011] [02] = 144'h 000000082212211020080884881041082000;  // FFFDB2D3BDD9680000 -0.2876820724517809 = 0.5 * ln( 1 + -1 * 2^(-2+1) + (-1^2+ 0^2) * 2^(-2*2) )   n =  2   d_n = -1 
assign X[4'b1011] [03] = 144'h 000000020208404204800808800420801000;  // FFFEEE8717DD800000 -0.1335313926245226 = 0.5 * ln( 1 + -1 * 2^(-3+1) + (-1^2+ 0^2) * 2^(-2*3) )   n =  3   d_n = -1 
assign X[4'b1011] [04] = 144'h 000000008020211210841112010812002040;  // FFFF7BD33A53100000 -0.0645385211375712 = 0.5 * ln( 1 + -1 * 2^(-4+1) + (-1^2+ 0^2) * 2^(-2*4) )   n =  4   d_n = -1 
assign X[4'b1011] [05] = 144'h 000000002002008440440880481202020200;  // FFFFBEFA89D8600000 -0.0317486983145803 = 0.5 * ln( 1 + -1 * 2^(-5+1) + (-1^2+ 0^2) * 2^(-2*5) )   n =  5   d_n = -1 
assign X[4'b1011] [06] = 144'h 000000000800200211121102088111008204;  // FFFFDFBF534ED80000 -0.0157483569681392 = 0.5 * ln( 1 + -1 * 2^(-6+1) + (-1^2+ 0^2) * 2^(-2*6) )   n =  6   d_n = -1 
assign X[4'b1011] [07] = 144'h 000000000200020008444044408204048102;  // FFFFEFEFEA8A780000 -0.0078431774610259 = 0.5 * ln( 1 + -1 * 2^(-7+1) + (-1^2+ 0^2) * 2^(-2*7) )   n =  7   d_n = -1 
assign X[4'b1011] [08] = 144'h 000000000080002000211112111020844848;  // FFFFF7FBFD53500000 -0.0039138993211363 = 0.5 * ln( 1 + -1 * 2^(-8+1) + (-1^2+ 0^2) * 2^(-2*8) )   n =  8   d_n = -1 
assign X[4'b1011] [09] = 144'h 000000000020000200008444404444080880;  // FFFFFBFEFFAA880000 -0.0019550348358034 = 0.5 * ln( 1 + -1 * 2^(-9+1) + (-1^2+ 0^2) * 2^(-2*9) )   n =  9   d_n = -1 
assign X[4'b1011] [10] = 144'h 000000000008000020000211111211110202;  // FFFFFDFFBFF5500000 -0.0009770396478266 = 0.5 * ln( 1 + -1 * 2^(-10+1) + (-1^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = -1 
assign X[4'b1011] [11] = 144'h 000000000002000002000008444440444440;  // FFFFFEFFEFFEA80000 -0.0004884004981089 = 0.5 * ln( 1 + -1 * 2^(-11+1) + (-1^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = -1 
assign X[4'b1011] [12] = 144'h 000000000000800000200000211111121111;  // FFFFFF7FFBFFD80000 -0.0002441704321739 = 0.5 * ln( 1 + -1 * 2^(-12+1) + (-1^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = -1 
assign X[4'b1011] [13] = 144'h 000000000000200000020000008444444044;  // FFFFFFBFFEFFF80000 -0.0001220777636870 = 0.5 * ln( 1 + -1 * 2^(-13+1) + (-1^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = -1 
assign X[4'b1011] [14] = 144'h 000000000000080000002000000211111110;  // FFFFFFDFFFC0000000 -0.0000610370189709 = 0.5 * ln( 1 + -1 * 2^(-14+1) + (-1^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = -1 
assign X[4'b1011] [15] = 144'h 000000000000020000000200000008444444;  // FFFFFFEFFFF0000000 -0.0000305180437958 = 0.5 * ln( 1 + -1 * 2^(-15+1) + (-1^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = -1 
assign X[4'b1011] [16] = 144'h 000000000000008000000020000000088888;  // FFFFFFF7FFFC000000 -0.0000152589054790 = 0.5 * ln( 1 + -1 * 2^(-16+1) + (-1^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = -1 
assign X[4'b1011] [17] = 144'h 000000000000002000000002000000002222;  // FFFFFFFBFFFF000000 -0.0000076294236352 = 0.5 * ln( 1 + -1 * 2^(-17+1) + (-1^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = -1 
assign X[4'b1011] [18] = 144'h 000000000000000800000000200000000088;  // FFFFFFFDFFFFC00000 -0.0000038147045416 = 0.5 * ln( 1 + -1 * 2^(-18+1) + (-1^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = -1 
assign X[4'b1011] [19] = 144'h 000000000000000200000000020000000002;  // FFFFFFFEFFFFF00000 -0.0000019073504518 = 0.5 * ln( 1 + -1 * 2^(-19+1) + (-1^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = -1 
assign X[4'b1011] [20] = 144'h 000000000000000080000000002000000000;  // FFFFFFFF7FFFF80000 -0.0000009536747712 = 0.5 * ln( 1 + -1 * 2^(-20+1) + (-1^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = -1 
assign X[4'b1011] [21] = 144'h 000000000000000020000000000200000000;  // FFFFFFFFC000000000 -0.0000004768372719 = 0.5 * ln( 1 + -1 * 2^(-21+1) + (-1^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = -1 
assign X[4'b1011] [22] = 144'h 000000000000000008000000000020000000;  // FFFFFFFFE000000000 -0.0000002384186075 = 0.5 * ln( 1 + -1 * 2^(-22+1) + (-1^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = -1 
assign X[4'b1011] [23] = 144'h 000000000000000002000000000002000000;  // FFFFFFFFF000000000 -0.0000001192092967 = 0.5 * ln( 1 + -1 * 2^(-23+1) + (-1^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = -1 
assign X[4'b1011] [24] = 144'h 000000000000000000800000000000200000;  // FFFFFFFFF800000000 -0.0000000596046466 = 0.5 * ln( 1 + -1 * 2^(-24+1) + (-1^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = -1 
assign X[4'b1011] [25] = 144'h 000000000000000000200000000000020000;  // FFFFFFFFFC00000000 -0.0000000298023228 = 0.5 * ln( 1 + -1 * 2^(-25+1) + (-1^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = -1 
assign X[4'b1011] [26] = 144'h 000000000000000000080000000000002000;  // FFFFFFFFFE00000000 -0.0000000149011613 = 0.5 * ln( 1 + -1 * 2^(-26+1) + (-1^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = -1 
assign X[4'b1011] [27] = 144'h 000000000000000000020000000000000200;  // FFFFFFFFFF00000000 -0.0000000074505806 = 0.5 * ln( 1 + -1 * 2^(-27+1) + (-1^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = -1 
assign X[4'b1011] [28] = 144'h 000000000000000000008000000000000020;  // FFFFFFFFFF80000000 -0.0000000037252903 = 0.5 * ln( 1 + -1 * 2^(-28+1) + (-1^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = -1 
assign X[4'b1011] [29] = 144'h 000000000000000000002000000000000002;  // FFFFFFFFFFC0000000 -0.0000000018626452 = 0.5 * ln( 1 + -1 * 2^(-29+1) + (-1^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = -1 
assign X[4'b1011] [30] = 144'h 000000000000000000000800000000000000;  // FFFFFFFFFFE0000000 -0.0000000009313226 = 0.5 * ln( 1 + -1 * 2^(-30+1) + (-1^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = -1 
assign X[4'b1011] [31] = 144'h 000000000000000000000200000000000000;  // FFFFFFFFFFF0000000 -0.0000000004656613 = 0.5 * ln( 1 + -1 * 2^(-31+1) + (-1^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = -1 
assign X[4'b1011] [32] = 144'h 000000000000000000000080000000000000;  // FFFFFFFFFFF8000000 -0.0000000002328306 = 0.5 * ln( 1 + -1 * 2^(-32+1) + (-1^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = -1 
assign X[4'b1011] [33] = 144'h 000000000000000000000020000000000000;  // FFFFFFFFFFFC000000 -0.0000000001164153 = 0.5 * ln( 1 + -1 * 2^(-33+1) + (-1^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = -1 
assign X[4'b1011] [34] = 144'h 000000000000000000000008000000000000;  // FFFFFFFFFFFE000000 -0.0000000000582077 = 0.5 * ln( 1 + -1 * 2^(-34+1) + (-1^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = -1 
assign X[4'b1011] [35] = 144'h 000000000000000000000002000000000000;  // FFFFFFFFFFFF000000 -0.0000000000291038 = 0.5 * ln( 1 + -1 * 2^(-35+1) + (-1^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = -1 
assign X[4'b1011] [36] = 144'h 000000000000000000000000800000000000;  // FFFFFFFFFFFF800000 -0.0000000000145519 = 0.5 * ln( 1 + -1 * 2^(-36+1) + (-1^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = -1 
assign X[4'b1011] [37] = 144'h 000000000000000000000000200000000000;  // FFFFFFFFFFFFC00000 -0.0000000000072760 = 0.5 * ln( 1 + -1 * 2^(-37+1) + (-1^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = -1 
assign X[4'b1011] [38] = 144'h 000000000000000000000000080000000000;  // FFFFFFFFFFFFE00000 -0.0000000000036380 = 0.5 * ln( 1 + -1 * 2^(-38+1) + (-1^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = -1 
assign X[4'b1011] [39] = 144'h 000000000000000000000000020000000000;  // FFFFFFFFFFFFF00000 -0.0000000000018190 = 0.5 * ln( 1 + -1 * 2^(-39+1) + (-1^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = -1 
assign X[4'b1011] [40] = 144'h 000000000000000000000000008000000000;  // FFFFFFFFFFFFF80000 -0.0000000000009095 = 0.5 * ln( 1 + -1 * 2^(-40+1) + (-1^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = -1 
assign X[4'b1011] [41] = 144'h 000000000000000000000000002000000000;  // FFFFFFFFFFFFF80000 -0.0000000000004547 = 0.5 * ln( 1 + -1 * 2^(-41+1) + (-1^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = -1 
assign X[4'b1011] [42] = 144'h 000000000000000000000000000800000000;  // 1000000000000000000 -0.0000000000002274 = 0.5 * ln( 1 + -1 * 2^(-42+1) + (-1^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = -1 
assign X[4'b1011] [43] = 144'h 000000000000000000000000000200000000;  // 1000000000000000000 -0.0000000000001137 = 0.5 * ln( 1 + -1 * 2^(-43+1) + (-1^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = -1 
assign X[4'b1011] [44] = 144'h 000000000000000000000000000080000000;  // 1000000000000000000 -0.0000000000000568 = 0.5 * ln( 1 + -1 * 2^(-44+1) + (-1^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = -1 
assign X[4'b1011] [45] = 144'h 000000000000000000000000000020000000;  // 1000000000000000000 -0.0000000000000284 = 0.5 * ln( 1 + -1 * 2^(-45+1) + (-1^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = -1 
assign X[4'b1011] [46] = 144'h 000000000000000000000000000008000000;  // 1000000000000000000 -0.0000000000000142 = 0.5 * ln( 1 + -1 * 2^(-46+1) + (-1^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = -1 
assign X[4'b1011] [47] = 144'h 000000000000000000000000000002000000;  // 1000000000000000000 -0.0000000000000071 = 0.5 * ln( 1 + -1 * 2^(-47+1) + (-1^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = -1 
assign X[4'b1011] [48] = 144'h 000000000000000000000000000000800000;  // 1000000000000000000 -0.0000000000000036 = 0.5 * ln( 1 + -1 * 2^(-48+1) + (-1^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = -1 
assign X[4'b1011] [49] = 144'h 000000000000000000000000000000200000;  // 1000000000000000000 -0.0000000000000018 = 0.5 * ln( 1 + -1 * 2^(-49+1) + (-1^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = -1 
assign X[4'b1011] [50] = 144'h 000000000000000000000000000000080000;  // 1000000000000000000 -0.0000000000000009 = 0.5 * ln( 1 + -1 * 2^(-50+1) + (-1^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = -1 
assign X[4'b1011] [51] = 144'h 000000000000000000000000000000020000;  // 1000000000000000000 -0.0000000000000004 = 0.5 * ln( 1 + -1 * 2^(-51+1) + (-1^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = -1 
assign X[4'b1011] [52] = 144'h 000000000000000000000000000000008000;  // 1000000000000000000 -0.0000000000000002 = 0.5 * ln( 1 + -1 * 2^(-52+1) + (-1^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = -1 
assign X[4'b1011] [53] = 144'h 000000000000000000000000000000002000;  // 1000000000000000000 -0.0000000000000001 = 0.5 * ln( 1 + -1 * 2^(-53+1) + (-1^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = -1 
assign X[4'b1011] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-54+1) + (-1^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = -1 
assign X[4'b1011] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-55+1) + (-1^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = -1 
assign X[4'b1011] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-56+1) + (-1^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = -1 
assign X[4'b1011] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-57+1) + (-1^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = -1 
assign X[4'b1011] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-58+1) + (-1^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = -1 
assign X[4'b1011] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-59+1) + (-1^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = -1 
assign X[4'b1011] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-60+1) + (-1^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = -1 
assign X[4'b1011] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-61+1) + (-1^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = -1 
assign X[4'b1011] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-62+1) + (-1^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = -1 
assign X[4'b1011] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-63+1) + (-1^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = -1 
assign X[4'b1011] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-64+1) + (-1^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = -1 
assign X[4'b1100] [01] = 144'h 000000010810400020081021211121010400;  // 0000E47FBE3CD4D128 +0.1115717756571049 = 0.5 * ln( 1 +  0 * 2^(-1+1) + ( 0^2+-1^2) * 2^(-2*1) )   n =  1   d_n = -0-1i 
assign X[4'b1100] [02] = 144'h 000000001008011048048000041220111100;  // 00003E14618022C552 +0.0303123109082174 = 0.5 * ln( 1 +  0 * 2^(-2+1) + ( 0^2+-1^2) * 2^(-2*2) )   n =  2   d_n = -0-1i 
assign X[4'b1100] [03] = 144'h 000000000100080011104880400800042120;  // 00000FE054587E01CC +0.0077520932679826 = 0.5 * ln( 1 +  0 * 2^(-3+1) + ( 0^2+-1^2) * 2^(-2*3) )   n =  3   d_n = -0-1i 
assign X[4'b1100] [04] = 144'h 000000000010000800011110488804048404;  // 000003FE01545621A1 +0.0019493202078287 = 0.5 * ln( 1 +  0 * 2^(-4+1) + ( 0^2+-1^2) * 2^(-2*4) )   n =  4   d_n = -0-1i 
assign X[4'b1100] [05] = 144'h 000000000001000008000011111048888084;  // 000000FFE00554557A +0.0004880429865277 = 0.5 * ln( 1 +  0 * 2^(-5+1) + ( 0^2+-1^2) * 2^(-2*5) )   n =  5   d_n = -0-1i 
assign X[4'b1100] [06] = 144'h 000000000000100000080000011111100448;  // 0000003FFE00155425 +0.0001220554137636 = 0.5 * ln( 1 +  0 * 2^(-6+1) + ( 0^2+-1^2) * 2^(-2*6) )   n =  6   d_n = -0-1i 
assign X[4'b1100] [07] = 144'h 000000000000010000000800000011111110;  // 0000000FFFE0005554 +0.0000305166468403 = 0.5 * ln( 1 +  0 * 2^(-7+1) + ( 0^2+-1^2) * 2^(-2*7) )   n =  7   d_n = -0-1i 
assign X[4'b1100] [08] = 144'h 000000000000001000000008000000011111;  // 00000003FFFE000155 +0.0000076293363242 = 0.5 * ln( 1 +  0 * 2^(-8+1) + ( 0^2+-1^2) * 2^(-2*8) )   n =  8   d_n = -0-1i 
assign X[4'b1100] [09] = 144'h 000000000000000100000000080000000012;  // 00000000FFFFE00003 +0.0000019073449948 = 0.5 * ln( 1 +  0 * 2^(-9+1) + ( 0^2+-1^2) * 2^(-2*9) )   n =  9   d_n = -0-1i 
assign X[4'b1100] [10] = 144'h 000000000000000010000000000800000000;  // 000000003FFFFE0000 +0.0000004768369308 = 0.5 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+-1^2) * 2^(-2*10) )   n = 10   d_n = -0-1i 
assign X[4'b1100] [11] = 144'h 000000000000000001000000000008000000;  // 000000000FFFFFE000 +0.0000001192092753 = 0.5 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+-1^2) * 2^(-2*11) )   n = 11   d_n = -0-1i 
assign X[4'b1100] [12] = 144'h 000000000000000000100000000000080000;  // 0000000003FFFFFE00 +0.0000000298023215 = 0.5 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+-1^2) * 2^(-2*12) )   n = 12   d_n = -0-1i 
assign X[4'b1100] [13] = 144'h 000000000000000000010000000000000200;  // 0000000000FFFFFFF0 +0.0000000074505806 = 0.5 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+-1^2) * 2^(-2*13) )   n = 13   d_n = -0-1i 
assign X[4'b1100] [14] = 144'h 000000000000000000001000000000000002;  // 00000000003FFFFFFF +0.0000000018626451 = 0.5 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+-1^2) * 2^(-2*14) )   n = 14   d_n = -0-1i 
assign X[4'b1100] [15] = 144'h 000000000000000000000100000000000000;  // 00000000000FFFFFFF +0.0000000004656613 = 0.5 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+-1^2) * 2^(-2*15) )   n = 15   d_n = -0-1i 
assign X[4'b1100] [16] = 144'h 000000000000000000000010000000000000;  // 000000000003FFFFFF +0.0000000001164153 = 0.5 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+-1^2) * 2^(-2*16) )   n = 16   d_n = -0-1i 
assign X[4'b1100] [17] = 144'h 000000000000000000000001000000000000;  // 000000000000FFFFFF +0.0000000000291038 = 0.5 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+-1^2) * 2^(-2*17) )   n = 17   d_n = -0-1i 
assign X[4'b1100] [18] = 144'h 000000000000000000000000100000000000;  // 0000000000003FFFFF +0.0000000000072760 = 0.5 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+-1^2) * 2^(-2*18) )   n = 18   d_n = -0-1i 
assign X[4'b1100] [19] = 144'h 000000000000000000000000010000000000;  // 0000000000000FFFFF +0.0000000000018190 = 0.5 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+-1^2) * 2^(-2*19) )   n = 19   d_n = -0-1i 
assign X[4'b1100] [20] = 144'h 000000000000000000000000001000000000;  // 00000000000003FFFF +0.0000000000004547 = 0.5 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+-1^2) * 2^(-2*20) )   n = 20   d_n = -0-1i 
assign X[4'b1100] [21] = 144'h 000000000000000000000000000100000000;  // 00000000000000FFFF +0.0000000000001137 = 0.5 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+-1^2) * 2^(-2*21) )   n = 21   d_n = -0-1i 
assign X[4'b1100] [22] = 144'h 000000000000000000000000000010000000;  // 000000000000003FFF +0.0000000000000284 = 0.5 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+-1^2) * 2^(-2*22) )   n = 22   d_n = -0-1i 
assign X[4'b1100] [23] = 144'h 000000000000000000000000000001000000;  // 000000000000000FFF +0.0000000000000071 = 0.5 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+-1^2) * 2^(-2*23) )   n = 23   d_n = -0-1i 
assign X[4'b1100] [24] = 144'h 000000000000000000000000000000100000;  // 0000000000000003FF +0.0000000000000018 = 0.5 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+-1^2) * 2^(-2*24) )   n = 24   d_n = -0-1i 
assign X[4'b1100] [25] = 144'h 000000000000000000000000000000010000;  // 0000000000000000FF +0.0000000000000004 = 0.5 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+-1^2) * 2^(-2*25) )   n = 25   d_n = -0-1i 
assign X[4'b1100] [26] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+-1^2) * 2^(-2*26) )   n = 26   d_n = -0-1i 
assign X[4'b1100] [27] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+-1^2) * 2^(-2*27) )   n = 27   d_n = -0-1i 
assign X[4'b1100] [28] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+-1^2) * 2^(-2*28) )   n = 28   d_n = -0-1i 
assign X[4'b1100] [29] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+-1^2) * 2^(-2*29) )   n = 29   d_n = -0-1i 
assign X[4'b1100] [30] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+-1^2) * 2^(-2*30) )   n = 30   d_n = -0-1i 
assign X[4'b1100] [31] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+-1^2) * 2^(-2*31) )   n = 31   d_n = -0-1i 
assign X[4'b1100] [32] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+-1^2) * 2^(-2*32) )   n = 32   d_n = -0-1i 
assign X[4'b1100] [33] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+-1^2) * 2^(-2*33) )   n = 33   d_n = -0-1i 
assign X[4'b1100] [34] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+-1^2) * 2^(-2*34) )   n = 34   d_n = -0-1i 
assign X[4'b1100] [35] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+-1^2) * 2^(-2*35) )   n = 35   d_n = -0-1i 
assign X[4'b1100] [36] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+-1^2) * 2^(-2*36) )   n = 36   d_n = -0-1i 
assign X[4'b1100] [37] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+-1^2) * 2^(-2*37) )   n = 37   d_n = -0-1i 
assign X[4'b1100] [38] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+-1^2) * 2^(-2*38) )   n = 38   d_n = -0-1i 
assign X[4'b1100] [39] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+-1^2) * 2^(-2*39) )   n = 39   d_n = -0-1i 
assign X[4'b1100] [40] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+-1^2) * 2^(-2*40) )   n = 40   d_n = -0-1i 
assign X[4'b1100] [41] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+-1^2) * 2^(-2*41) )   n = 41   d_n = -0-1i 
assign X[4'b1100] [42] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+-1^2) * 2^(-2*42) )   n = 42   d_n = -0-1i 
assign X[4'b1100] [43] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+-1^2) * 2^(-2*43) )   n = 43   d_n = -0-1i 
assign X[4'b1100] [44] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+-1^2) * 2^(-2*44) )   n = 44   d_n = -0-1i 
assign X[4'b1100] [45] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+-1^2) * 2^(-2*45) )   n = 45   d_n = -0-1i 
assign X[4'b1100] [46] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+-1^2) * 2^(-2*46) )   n = 46   d_n = -0-1i 
assign X[4'b1100] [47] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+-1^2) * 2^(-2*47) )   n = 47   d_n = -0-1i 
assign X[4'b1100] [48] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+-1^2) * 2^(-2*48) )   n = 48   d_n = -0-1i 
assign X[4'b1100] [49] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+-1^2) * 2^(-2*49) )   n = 49   d_n = -0-1i 
assign X[4'b1100] [50] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+-1^2) * 2^(-2*50) )   n = 50   d_n = -0-1i 
assign X[4'b1100] [51] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+-1^2) * 2^(-2*51) )   n = 51   d_n = -0-1i 
assign X[4'b1100] [52] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+-1^2) * 2^(-2*52) )   n = 52   d_n = -0-1i 
assign X[4'b1100] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+-1^2) * 2^(-2*53) )   n = 53   d_n = -0-1i 
assign X[4'b1100] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+-1^2) * 2^(-2*54) )   n = 54   d_n = -0-1i 
assign X[4'b1100] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+-1^2) * 2^(-2*55) )   n = 55   d_n = -0-1i 
assign X[4'b1100] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+-1^2) * 2^(-2*56) )   n = 56   d_n = -0-1i 
assign X[4'b1100] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+-1^2) * 2^(-2*57) )   n = 57   d_n = -0-1i 
assign X[4'b1100] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+-1^2) * 2^(-2*58) )   n = 58   d_n = -0-1i 
assign X[4'b1100] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+-1^2) * 2^(-2*59) )   n = 59   d_n = -0-1i 
assign X[4'b1100] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+-1^2) * 2^(-2*60) )   n = 60   d_n = -0-1i 
assign X[4'b1100] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+-1^2) * 2^(-2*61) )   n = 61   d_n = -0-1i 
assign X[4'b1100] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+-1^2) * 2^(-2*62) )   n = 62   d_n = -0-1i 
assign X[4'b1100] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+-1^2) * 2^(-2*63) )   n = 63   d_n = -0-1i 
assign X[4'b1100] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+-1^2) * 2^(-2*64) )   n = 64   d_n = -0-1i 
assign X[4'b1101] [01] = 144'h 000000108444104004080420042001020000;  // 0003AA481E1C1C0F20 +0.4581453659370776 = 0.5 * ln( 1 +  1 * 2^(-1+1) + ( 1^2+-1^2) * 2^(-2*1) )   n =  1   d_n = 1-1i 
assign X[4'b1101] [02] = 144'h 000000040201044100880022020042084400;  // 0001F128F5FAF06EA0 +0.2427539078908503 = 0.5 * ln( 1 +  1 * 2^(-2+1) + ( 1^2+-1^2) * 2^(-2*2) )   n =  2   d_n = 1-1i 
assign X[4'b1101] [03] = 144'h 000000010008204120108222020402048000;  // 0000FDC8C36AF1F180 +0.1239180819522907 = 0.5 * ln( 1 +  1 * 2^(-3+1) + ( 1^2+-1^2) * 2^(-2*3) )   n =  3   d_n = 1-1i 
assign X[4'b1101] [04] = 144'h 000000004000220410112040820022220420;  // 00007FB244C76FAB1C +0.0623517392504787 = 0.5 * ln( 1 +  1 * 2^(-4+1) + ( 1^2+-1^2) * 2^(-2*4) )   n =  4   d_n = 1-1i 
assign X[4'b1101] [05] = 144'h 000000001000008821040412108204480088;  // 00003FF5D2233725F6 +0.0312305848118681 = 0.5 * ln( 1 +  1 * 2^(-5+1) + ( 1^2+-1^2) * 2^(-2*5) )   n =  5   d_n = 1-1i 
assign X[4'b1101] [06] = 144'h 000000000400000222044101011210441080;  // 00001FFEB291134A38 +0.0156225157283291 = 0.5 * ln( 1 +  1 * 2^(-6+1) + ( 1^2+-1^2) * 2^(-2*6) )   n =  6   d_n = 1-1i 
assign X[4'b1101] [07] = 144'h 000000000100000008882110404041212102;  // 00000FFFD5D4888CCF +0.0078121858105703 = 0.5 * ln( 1 +  1 * 2^(-7+1) + ( 1^2+-1^2) * 2^(-2*7) )   n =  7   d_n = 1-1i 
assign X[4'b1101] [08] = 144'h 000000000040000000222204441010101044;  // 000007FFFAB2A4444A +0.0039062104956732 = 0.5 * ln( 1 +  1 * 2^(-8+1) + ( 1^2+-1^2) * 2^(-2*8) )   n =  8   d_n = 1-1i 
assign X[4'b1101] [09] = 144'h 000000000010000000008888211104040440;  // 000003FFFF55D52228 +0.0019531200474755 = 0.5 * ln( 1 +  1 * 2^(-9+1) + ( 1^2+-1^2) * 2^(-2*9) )   n =  9   d_n = 1-1i 
assign X[4'b1101] [10] = 144'h 000000000004000000000222220444412101;  // 000001FFFFEAB2A8D1 +0.0009765618800270 = 0.5 * ln( 1 +  1 * 2^(-10+1) + ( 1^2+-1^2) * 2^(-2*10) )   n = 10   d_n = 1-1i 
assign X[4'b1101] [11] = 144'h 000000000001000000000008888821111044;  // 000000FFFFFD55D54A +0.0004882811724466 = 0.5 * ln( 1 +  1 * 2^(-11+1) + ( 1^2+-1^2) * 2^(-2*11) )   n = 11   d_n = 1-1i 
assign X[4'b1101] [12] = 144'h 000000000000400000000000222222044444;  // 0000007FFFFFAAB2AA +0.0002441406153023 = 0.5 * ln( 1 +  1 * 2^(-12+1) + ( 1^2+-1^2) * 2^(-2*12) )   n = 12   d_n = 1-1i 
assign X[4'b1101] [13] = 144'h 000000000000100000000000008888888411;  // 0000003FFFFFF555A5 +0.0001220703112875 = 0.5 * ln( 1 +  1 * 2^(-13+1) + ( 1^2+-1^2) * 2^(-2*13) )   n = 13   d_n = 1-1i 
assign X[4'b1101] [14] = 144'h 000000000000040000000000000222222200;  // 0000001FFFFFFEAAAF +0.0000610351560984 = 0.5 * ln( 1 +  1 * 2^(-14+1) + ( 1^2+-1^2) * 2^(-2*14) )   n = 14   d_n = 1-1i 
assign X[4'b1101] [15] = 144'h 000000000000010000000000000008888888;  // 0000000FFFFFFFD555 +0.0000305175781061 = 0.5 * ln( 1 +  1 * 2^(-15+1) + ( 1^2+-1^2) * 2^(-2*15) )   n = 15   d_n = 1-1i 
assign X[4'b1101] [16] = 144'h 000000000000004000000000000000844444;  // 00000007FFFFFFFAAA +0.0000152587890601 = 0.5 * ln( 1 +  1 * 2^(-16+1) + ( 1^2+-1^2) * 2^(-2*16) )   n = 16   d_n = 1-1i 
assign X[4'b1101] [17] = 144'h 000000000000001000000000000000021111;  // 00000003FFFFFFFF55 +0.0000076293945310 = 0.5 * ln( 1 +  1 * 2^(-17+1) + ( 1^2+-1^2) * 2^(-2*17) )   n = 17   d_n = 1-1i 
assign X[4'b1101] [18] = 144'h 000000000000000400000000000000000084;  // 00000001FFFFFFFFFA +0.0000038146972656 = 0.5 * ln( 1 +  1 * 2^(-18+1) + ( 1^2+-1^2) * 2^(-2*18) )   n = 18   d_n = 1-1i 
assign X[4'b1101] [19] = 144'h 000000000000000100000000000000000002;  // 00000000FFFFFFFFFF +0.0000019073486328 = 0.5 * ln( 1 +  1 * 2^(-19+1) + ( 1^2+-1^2) * 2^(-2*19) )   n = 19   d_n = 1-1i 
assign X[4'b1101] [20] = 144'h 000000000000000040000000000000000000;  // 000000007FFFFFFFFF +0.0000009536743164 = 0.5 * ln( 1 +  1 * 2^(-20+1) + ( 1^2+-1^2) * 2^(-2*20) )   n = 20   d_n = 1-1i 
assign X[4'b1101] [21] = 144'h 000000000000000010000000000000000000;  // 000000003FFFFFFFFF +0.0000004768371582 = 0.5 * ln( 1 +  1 * 2^(-21+1) + ( 1^2+-1^2) * 2^(-2*21) )   n = 21   d_n = 1-1i 
assign X[4'b1101] [22] = 144'h 000000000000000004000000000000000000;  // 000000001FFFFFFFFF +0.0000002384185791 = 0.5 * ln( 1 +  1 * 2^(-22+1) + ( 1^2+-1^2) * 2^(-2*22) )   n = 22   d_n = 1-1i 
assign X[4'b1101] [23] = 144'h 000000000000000001000000000000000000;  // 000000000FFFFFFFFF +0.0000001192092896 = 0.5 * ln( 1 +  1 * 2^(-23+1) + ( 1^2+-1^2) * 2^(-2*23) )   n = 23   d_n = 1-1i 
assign X[4'b1101] [24] = 144'h 000000000000000000400000000000000000;  // 0000000007FFFFFFFF +0.0000000596046448 = 0.5 * ln( 1 +  1 * 2^(-24+1) + ( 1^2+-1^2) * 2^(-2*24) )   n = 24   d_n = 1-1i 
assign X[4'b1101] [25] = 144'h 000000000000000000100000000000000000;  // 0000000003FFFFFFFF +0.0000000298023224 = 0.5 * ln( 1 +  1 * 2^(-25+1) + ( 1^2+-1^2) * 2^(-2*25) )   n = 25   d_n = 1-1i 
assign X[4'b1101] [26] = 144'h 000000000000000000040000000000002000;  // 0000000001FFFFFFC0 +0.0000000149011611 = 0.5 * ln( 1 +  1 * 2^(-26+1) + ( 1^2+-1^2) * 2^(-2*26) )   n = 26   d_n = 1-1i 
assign X[4'b1101] [27] = 144'h 000000000000000000010000000000000200;  // 0000000000FFFFFFF0 +0.0000000074505806 = 0.5 * ln( 1 +  1 * 2^(-27+1) + ( 1^2+-1^2) * 2^(-2*27) )   n = 27   d_n = 1-1i 
assign X[4'b1101] [28] = 144'h 000000000000000000004000000000000020;  // 00000000007FFFFFFC +0.0000000037252903 = 0.5 * ln( 1 +  1 * 2^(-28+1) + ( 1^2+-1^2) * 2^(-2*28) )   n = 28   d_n = 1-1i 
assign X[4'b1101] [29] = 144'h 000000000000000000001000000000000002;  // 00000000003FFFFFFF +0.0000000018626451 = 0.5 * ln( 1 +  1 * 2^(-29+1) + ( 1^2+-1^2) * 2^(-2*29) )   n = 29   d_n = 1-1i 
assign X[4'b1101] [30] = 144'h 000000000000000000000400000000000000;  // 00000000001FFFFFFF +0.0000000009313226 = 0.5 * ln( 1 +  1 * 2^(-30+1) + ( 1^2+-1^2) * 2^(-2*30) )   n = 30   d_n = 1-1i 
assign X[4'b1101] [31] = 144'h 000000000000000000000100000000000000;  // 00000000000FFFFFFF +0.0000000004656613 = 0.5 * ln( 1 +  1 * 2^(-31+1) + ( 1^2+-1^2) * 2^(-2*31) )   n = 31   d_n = 1-1i 
assign X[4'b1101] [32] = 144'h 000000000000000000000040000000000000;  // 000000000007FFFFFF +0.0000000002328306 = 0.5 * ln( 1 +  1 * 2^(-32+1) + ( 1^2+-1^2) * 2^(-2*32) )   n = 32   d_n = 1-1i 
assign X[4'b1101] [33] = 144'h 000000000000000000000010000000000000;  // 000000000003FFFFFF +0.0000000001164153 = 0.5 * ln( 1 +  1 * 2^(-33+1) + ( 1^2+-1^2) * 2^(-2*33) )   n = 33   d_n = 1-1i 
assign X[4'b1101] [34] = 144'h 000000000000000000000004000000000000;  // 000000000001FFFFFF +0.0000000000582077 = 0.5 * ln( 1 +  1 * 2^(-34+1) + ( 1^2+-1^2) * 2^(-2*34) )   n = 34   d_n = 1-1i 
assign X[4'b1101] [35] = 144'h 000000000000000000000001000000000000;  // 000000000000FFFFFF +0.0000000000291038 = 0.5 * ln( 1 +  1 * 2^(-35+1) + ( 1^2+-1^2) * 2^(-2*35) )   n = 35   d_n = 1-1i 
assign X[4'b1101] [36] = 144'h 000000000000000000000000400000000000;  // 0000000000007FFFFF +0.0000000000145519 = 0.5 * ln( 1 +  1 * 2^(-36+1) + ( 1^2+-1^2) * 2^(-2*36) )   n = 36   d_n = 1-1i 
assign X[4'b1101] [37] = 144'h 000000000000000000000000100000000000;  // 0000000000003FFFFF +0.0000000000072760 = 0.5 * ln( 1 +  1 * 2^(-37+1) + ( 1^2+-1^2) * 2^(-2*37) )   n = 37   d_n = 1-1i 
assign X[4'b1101] [38] = 144'h 000000000000000000000000040000000000;  // 0000000000001FFFFF +0.0000000000036380 = 0.5 * ln( 1 +  1 * 2^(-38+1) + ( 1^2+-1^2) * 2^(-2*38) )   n = 38   d_n = 1-1i 
assign X[4'b1101] [39] = 144'h 000000000000000000000000010000000000;  // 0000000000000FFFFF +0.0000000000018190 = 0.5 * ln( 1 +  1 * 2^(-39+1) + ( 1^2+-1^2) * 2^(-2*39) )   n = 39   d_n = 1-1i 
assign X[4'b1101] [40] = 144'h 000000000000000000000000004000000000;  // 00000000000007FFFF +0.0000000000009095 = 0.5 * ln( 1 +  1 * 2^(-40+1) + ( 1^2+-1^2) * 2^(-2*40) )   n = 40   d_n = 1-1i 
assign X[4'b1101] [41] = 144'h 000000000000000000000000001000000000;  // 00000000000003FFFF +0.0000000000004547 = 0.5 * ln( 1 +  1 * 2^(-41+1) + ( 1^2+-1^2) * 2^(-2*41) )   n = 41   d_n = 1-1i 
assign X[4'b1101] [42] = 144'h 000000000000000000000000000400000000;  // 00000000000001FFFF +0.0000000000002274 = 0.5 * ln( 1 +  1 * 2^(-42+1) + ( 1^2+-1^2) * 2^(-2*42) )   n = 42   d_n = 1-1i 
assign X[4'b1101] [43] = 144'h 000000000000000000000000000100000000;  // 00000000000000FFFF +0.0000000000001137 = 0.5 * ln( 1 +  1 * 2^(-43+1) + ( 1^2+-1^2) * 2^(-2*43) )   n = 43   d_n = 1-1i 
assign X[4'b1101] [44] = 144'h 000000000000000000000000000040000000;  // 000000000000007FFF +0.0000000000000568 = 0.5 * ln( 1 +  1 * 2^(-44+1) + ( 1^2+-1^2) * 2^(-2*44) )   n = 44   d_n = 1-1i 
assign X[4'b1101] [45] = 144'h 000000000000000000000000000010000000;  // 000000000000003FFF +0.0000000000000284 = 0.5 * ln( 1 +  1 * 2^(-45+1) + ( 1^2+-1^2) * 2^(-2*45) )   n = 45   d_n = 1-1i 
assign X[4'b1101] [46] = 144'h 000000000000000000000000000004000000;  // 000000000000001FFF +0.0000000000000142 = 0.5 * ln( 1 +  1 * 2^(-46+1) + ( 1^2+-1^2) * 2^(-2*46) )   n = 46   d_n = 1-1i 
assign X[4'b1101] [47] = 144'h 000000000000000000000000000001000000;  // 000000000000000FFF +0.0000000000000071 = 0.5 * ln( 1 +  1 * 2^(-47+1) + ( 1^2+-1^2) * 2^(-2*47) )   n = 47   d_n = 1-1i 
assign X[4'b1101] [48] = 144'h 000000000000000000000000000000400000;  // 0000000000000007FF +0.0000000000000036 = 0.5 * ln( 1 +  1 * 2^(-48+1) + ( 1^2+-1^2) * 2^(-2*48) )   n = 48   d_n = 1-1i 
assign X[4'b1101] [49] = 144'h 000000000000000000000000000000100000;  // 0000000000000003FF +0.0000000000000018 = 0.5 * ln( 1 +  1 * 2^(-49+1) + ( 1^2+-1^2) * 2^(-2*49) )   n = 49   d_n = 1-1i 
assign X[4'b1101] [50] = 144'h 000000000000000000000000000000040000;  // 0000000000000001FF +0.0000000000000009 = 0.5 * ln( 1 +  1 * 2^(-50+1) + ( 1^2+-1^2) * 2^(-2*50) )   n = 50   d_n = 1-1i 
assign X[4'b1101] [51] = 144'h 000000000000000000000000000000010000;  // 0000000000000000FF +0.0000000000000004 = 0.5 * ln( 1 +  1 * 2^(-51+1) + ( 1^2+-1^2) * 2^(-2*51) )   n = 51   d_n = 1-1i 
assign X[4'b1101] [52] = 144'h 000000000000000000000000000000004000;  // 00000000000000007F +0.0000000000000002 = 0.5 * ln( 1 +  1 * 2^(-52+1) + ( 1^2+-1^2) * 2^(-2*52) )   n = 52   d_n = 1-1i 
assign X[4'b1101] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-53+1) + ( 1^2+-1^2) * 2^(-2*53) )   n = 53   d_n = 1-1i 
assign X[4'b1101] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-54+1) + ( 1^2+-1^2) * 2^(-2*54) )   n = 54   d_n = 1-1i 
assign X[4'b1101] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-55+1) + ( 1^2+-1^2) * 2^(-2*55) )   n = 55   d_n = 1-1i 
assign X[4'b1101] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-56+1) + ( 1^2+-1^2) * 2^(-2*56) )   n = 56   d_n = 1-1i 
assign X[4'b1101] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-57+1) + ( 1^2+-1^2) * 2^(-2*57) )   n = 57   d_n = 1-1i 
assign X[4'b1101] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-58+1) + ( 1^2+-1^2) * 2^(-2*58) )   n = 58   d_n = 1-1i 
assign X[4'b1101] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-59+1) + ( 1^2+-1^2) * 2^(-2*59) )   n = 59   d_n = 1-1i 
assign X[4'b1101] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-60+1) + ( 1^2+-1^2) * 2^(-2*60) )   n = 60   d_n = 1-1i 
assign X[4'b1101] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-61+1) + ( 1^2+-1^2) * 2^(-2*61) )   n = 61   d_n = 1-1i 
assign X[4'b1101] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-62+1) + ( 1^2+-1^2) * 2^(-2*62) )   n = 62   d_n = 1-1i 
assign X[4'b1101] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-63+1) + ( 1^2+-1^2) * 2^(-2*63) )   n = 63   d_n = 1-1i 
assign X[4'b1101] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  1 * 2^(-64+1) + ( 1^2+-1^2) * 2^(-2*64) )   n = 64   d_n = 1-1i 
assign X[4'b1110] [01] = 144'h 000000010810400020081021211121010400;  // 0000E47FBE3CD4D128 +0.1115717756571049 = 0.5 * ln( 1 +  0 * 2^(-1+1) + ( 0^2+-1^2) * 2^(-2*1) )   n =  1   d_n = -0-1i 
assign X[4'b1110] [02] = 144'h 000000001008011048048000041220111100;  // 00003E14618022C552 +0.0303123109082174 = 0.5 * ln( 1 +  0 * 2^(-2+1) + ( 0^2+-1^2) * 2^(-2*2) )   n =  2   d_n = -0-1i 
assign X[4'b1110] [03] = 144'h 000000000100080011104880400800042120;  // 00000FE054587E01CC +0.0077520932679826 = 0.5 * ln( 1 +  0 * 2^(-3+1) + ( 0^2+-1^2) * 2^(-2*3) )   n =  3   d_n = -0-1i 
assign X[4'b1110] [04] = 144'h 000000000010000800011110488804048404;  // 000003FE01545621A1 +0.0019493202078287 = 0.5 * ln( 1 +  0 * 2^(-4+1) + ( 0^2+-1^2) * 2^(-2*4) )   n =  4   d_n = -0-1i 
assign X[4'b1110] [05] = 144'h 000000000001000008000011111048888084;  // 000000FFE00554557A +0.0004880429865277 = 0.5 * ln( 1 +  0 * 2^(-5+1) + ( 0^2+-1^2) * 2^(-2*5) )   n =  5   d_n = -0-1i 
assign X[4'b1110] [06] = 144'h 000000000000100000080000011111100448;  // 0000003FFE00155425 +0.0001220554137636 = 0.5 * ln( 1 +  0 * 2^(-6+1) + ( 0^2+-1^2) * 2^(-2*6) )   n =  6   d_n = -0-1i 
assign X[4'b1110] [07] = 144'h 000000000000010000000800000011111110;  // 0000000FFFE0005554 +0.0000305166468403 = 0.5 * ln( 1 +  0 * 2^(-7+1) + ( 0^2+-1^2) * 2^(-2*7) )   n =  7   d_n = -0-1i 
assign X[4'b1110] [08] = 144'h 000000000000001000000008000000011111;  // 00000003FFFE000155 +0.0000076293363242 = 0.5 * ln( 1 +  0 * 2^(-8+1) + ( 0^2+-1^2) * 2^(-2*8) )   n =  8   d_n = -0-1i 
assign X[4'b1110] [09] = 144'h 000000000000000100000000080000000012;  // 00000000FFFFE00003 +0.0000019073449948 = 0.5 * ln( 1 +  0 * 2^(-9+1) + ( 0^2+-1^2) * 2^(-2*9) )   n =  9   d_n = -0-1i 
assign X[4'b1110] [10] = 144'h 000000000000000010000000000800000000;  // 000000003FFFFE0000 +0.0000004768369308 = 0.5 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+-1^2) * 2^(-2*10) )   n = 10   d_n = -0-1i 
assign X[4'b1110] [11] = 144'h 000000000000000001000000000008000000;  // 000000000FFFFFE000 +0.0000001192092753 = 0.5 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+-1^2) * 2^(-2*11) )   n = 11   d_n = -0-1i 
assign X[4'b1110] [12] = 144'h 000000000000000000100000000000080000;  // 0000000003FFFFFE00 +0.0000000298023215 = 0.5 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+-1^2) * 2^(-2*12) )   n = 12   d_n = -0-1i 
assign X[4'b1110] [13] = 144'h 000000000000000000010000000000000200;  // 0000000000FFFFFFF0 +0.0000000074505806 = 0.5 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+-1^2) * 2^(-2*13) )   n = 13   d_n = -0-1i 
assign X[4'b1110] [14] = 144'h 000000000000000000001000000000000002;  // 00000000003FFFFFFF +0.0000000018626451 = 0.5 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+-1^2) * 2^(-2*14) )   n = 14   d_n = -0-1i 
assign X[4'b1110] [15] = 144'h 000000000000000000000100000000000000;  // 00000000000FFFFFFF +0.0000000004656613 = 0.5 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+-1^2) * 2^(-2*15) )   n = 15   d_n = -0-1i 
assign X[4'b1110] [16] = 144'h 000000000000000000000010000000000000;  // 000000000003FFFFFF +0.0000000001164153 = 0.5 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+-1^2) * 2^(-2*16) )   n = 16   d_n = -0-1i 
assign X[4'b1110] [17] = 144'h 000000000000000000000001000000000000;  // 000000000000FFFFFF +0.0000000000291038 = 0.5 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+-1^2) * 2^(-2*17) )   n = 17   d_n = -0-1i 
assign X[4'b1110] [18] = 144'h 000000000000000000000000100000000000;  // 0000000000003FFFFF +0.0000000000072760 = 0.5 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+-1^2) * 2^(-2*18) )   n = 18   d_n = -0-1i 
assign X[4'b1110] [19] = 144'h 000000000000000000000000010000000000;  // 0000000000000FFFFF +0.0000000000018190 = 0.5 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+-1^2) * 2^(-2*19) )   n = 19   d_n = -0-1i 
assign X[4'b1110] [20] = 144'h 000000000000000000000000001000000000;  // 00000000000003FFFF +0.0000000000004547 = 0.5 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+-1^2) * 2^(-2*20) )   n = 20   d_n = -0-1i 
assign X[4'b1110] [21] = 144'h 000000000000000000000000000100000000;  // 00000000000000FFFF +0.0000000000001137 = 0.5 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+-1^2) * 2^(-2*21) )   n = 21   d_n = -0-1i 
assign X[4'b1110] [22] = 144'h 000000000000000000000000000010000000;  // 000000000000003FFF +0.0000000000000284 = 0.5 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+-1^2) * 2^(-2*22) )   n = 22   d_n = -0-1i 
assign X[4'b1110] [23] = 144'h 000000000000000000000000000001000000;  // 000000000000000FFF +0.0000000000000071 = 0.5 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+-1^2) * 2^(-2*23) )   n = 23   d_n = -0-1i 
assign X[4'b1110] [24] = 144'h 000000000000000000000000000000100000;  // 0000000000000003FF +0.0000000000000018 = 0.5 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+-1^2) * 2^(-2*24) )   n = 24   d_n = -0-1i 
assign X[4'b1110] [25] = 144'h 000000000000000000000000000000010000;  // 0000000000000000FF +0.0000000000000004 = 0.5 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+-1^2) * 2^(-2*25) )   n = 25   d_n = -0-1i 
assign X[4'b1110] [26] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+-1^2) * 2^(-2*26) )   n = 26   d_n = -0-1i 
assign X[4'b1110] [27] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+-1^2) * 2^(-2*27) )   n = 27   d_n = -0-1i 
assign X[4'b1110] [28] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+-1^2) * 2^(-2*28) )   n = 28   d_n = -0-1i 
assign X[4'b1110] [29] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+-1^2) * 2^(-2*29) )   n = 29   d_n = -0-1i 
assign X[4'b1110] [30] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+-1^2) * 2^(-2*30) )   n = 30   d_n = -0-1i 
assign X[4'b1110] [31] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+-1^2) * 2^(-2*31) )   n = 31   d_n = -0-1i 
assign X[4'b1110] [32] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+-1^2) * 2^(-2*32) )   n = 32   d_n = -0-1i 
assign X[4'b1110] [33] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+-1^2) * 2^(-2*33) )   n = 33   d_n = -0-1i 
assign X[4'b1110] [34] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+-1^2) * 2^(-2*34) )   n = 34   d_n = -0-1i 
assign X[4'b1110] [35] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+-1^2) * 2^(-2*35) )   n = 35   d_n = -0-1i 
assign X[4'b1110] [36] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+-1^2) * 2^(-2*36) )   n = 36   d_n = -0-1i 
assign X[4'b1110] [37] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+-1^2) * 2^(-2*37) )   n = 37   d_n = -0-1i 
assign X[4'b1110] [38] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+-1^2) * 2^(-2*38) )   n = 38   d_n = -0-1i 
assign X[4'b1110] [39] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+-1^2) * 2^(-2*39) )   n = 39   d_n = -0-1i 
assign X[4'b1110] [40] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+-1^2) * 2^(-2*40) )   n = 40   d_n = -0-1i 
assign X[4'b1110] [41] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+-1^2) * 2^(-2*41) )   n = 41   d_n = -0-1i 
assign X[4'b1110] [42] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+-1^2) * 2^(-2*42) )   n = 42   d_n = -0-1i 
assign X[4'b1110] [43] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+-1^2) * 2^(-2*43) )   n = 43   d_n = -0-1i 
assign X[4'b1110] [44] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+-1^2) * 2^(-2*44) )   n = 44   d_n = -0-1i 
assign X[4'b1110] [45] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+-1^2) * 2^(-2*45) )   n = 45   d_n = -0-1i 
assign X[4'b1110] [46] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+-1^2) * 2^(-2*46) )   n = 46   d_n = -0-1i 
assign X[4'b1110] [47] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+-1^2) * 2^(-2*47) )   n = 47   d_n = -0-1i 
assign X[4'b1110] [48] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+-1^2) * 2^(-2*48) )   n = 48   d_n = -0-1i 
assign X[4'b1110] [49] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+-1^2) * 2^(-2*49) )   n = 49   d_n = -0-1i 
assign X[4'b1110] [50] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+-1^2) * 2^(-2*50) )   n = 50   d_n = -0-1i 
assign X[4'b1110] [51] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+-1^2) * 2^(-2*51) )   n = 51   d_n = -0-1i 
assign X[4'b1110] [52] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+-1^2) * 2^(-2*52) )   n = 52   d_n = -0-1i 
assign X[4'b1110] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+-1^2) * 2^(-2*53) )   n = 53   d_n = -0-1i 
assign X[4'b1110] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+-1^2) * 2^(-2*54) )   n = 54   d_n = -0-1i 
assign X[4'b1110] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+-1^2) * 2^(-2*55) )   n = 55   d_n = -0-1i 
assign X[4'b1110] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+-1^2) * 2^(-2*56) )   n = 56   d_n = -0-1i 
assign X[4'b1110] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+-1^2) * 2^(-2*57) )   n = 57   d_n = -0-1i 
assign X[4'b1110] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+-1^2) * 2^(-2*58) )   n = 58   d_n = -0-1i 
assign X[4'b1110] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+-1^2) * 2^(-2*59) )   n = 59   d_n = -0-1i 
assign X[4'b1110] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+-1^2) * 2^(-2*60) )   n = 60   d_n = -0-1i 
assign X[4'b1110] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+-1^2) * 2^(-2*61) )   n = 61   d_n = -0-1i 
assign X[4'b1110] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+-1^2) * 2^(-2*62) )   n = 62   d_n = -0-1i 
assign X[4'b1110] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+-1^2) * 2^(-2*63) )   n = 63   d_n = -0-1i 
assign X[4'b1110] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+-1^2) * 2^(-2*64) )   n = 64   d_n = -0-1i 
assign X[4'b1111] [01] = 144'h 000000211084108084000401208120041000;  // FFFD3A37A020B80000 -0.3465735902799726 = 0.5 * ln( 1 + -1 * 2^(-1+1) + (-1^2+-1^2) * 2^(-2*1) )   n =  1   d_n = -1-1i 
assign X[4'b1111] [02] = 144'h 000000080402208088084808810881121100;  // FFFE1EB75E5D900000 -0.2350018146228677 = 0.5 * ln( 1 + -1 * 2^(-2+1) + (-1^2+-1^2) * 2^(-2*2) )   n =  2   d_n = -1-1i 
assign X[4'b1111] [03] = 144'h 000000020012108204204484480448101040;  // FFFF03371C9A600000 -0.1234300389657629 = 0.5 * ln( 1 + -1 * 2^(-3+1) + (-1^2+-1^2) * 2^(-2*3) )   n =  3   d_n = -1-1i 
assign X[4'b1111] [04] = 144'h 000000008000480820220480410044444810;  // FFFF805DBB18900000 -0.0623212226036383 = 0.5 * ln( 1 + -1 * 2^(-4+1) + (-1^2+-1^2) * 2^(-2*4) )   n =  4   d_n = -1-1i 
assign X[4'b1111] [05] = 144'h 000000002000012212080820444108840110;  // FFFFC00B2DDCA80000 -0.0312286774668733 = 0.5 * ln( 1 + -1 * 2^(-5+1) + (-1^2+-1^2) * 2^(-2*5) )   n =  5   d_n = -1-1i 
assign X[4'b1111] [06] = 144'h 000000000800000488088202022044888440;  // FFFFE0015D6EF00000 -0.0156223965190538 = 0.5 * ln( 1 + -1 * 2^(-6+1) + (-1^2+-1^2) * 2^(-2*6) )   n =  6   d_n = -1-1i 
assign X[4'b1111] [07] = 144'h 000000000200000012221220808082120881;  // FFFFF0002B2B780000 -0.0078121783599899 = 0.5 * ln( 1 + -1 * 2^(-7+1) + (-1^2+-1^2) * 2^(-2*7) )   n =  7   d_n = -1-1i 
assign X[4'b1111] [08] = 144'h 000000000080000000488808882020202088;  // FFFFF800055D580000 -0.0039062100300119 = 0.5 * ln( 1 + -1 * 2^(-8+1) + (-1^2+-1^2) * 2^(-2*8) )   n =  8   d_n = -1-1i 
assign X[4'b1111] [09] = 144'h 000000000020000000012222122208080810;  // FFFFFC0000AB280000 -0.0019531200183716 = 0.5 * ln( 1 + -1 * 2^(-9+1) + (-1^2+-1^2) * 2^(-2*9) )   n =  9   d_n = -1-1i 
assign X[4'b1111] [10] = 144'h 000000000008000000000488880888820202;  // FFFFFE000015600000 -0.0009765618782081 = 0.5 * ln( 1 + -1 * 2^(-10+1) + (-1^2+-1^2) * 2^(-2*10) )   n = 10   d_n = -1-1i 
assign X[4'b1111] [11] = 144'h 000000000002000000000012222212222088;  // FFFFFF000002A80000 -0.0004882811723329 = 0.5 * ln( 1 + -1 * 2^(-11+1) + (-1^2+-1^2) * 2^(-2*11) )   n = 11   d_n = -1-1i 
assign X[4'b1111] [12] = 144'h 000000000000800000000000488888088888;  // FFFFFF800000580000 -0.0002441406152952 = 0.5 * ln( 1 + -1 * 2^(-12+1) + (-1^2+-1^2) * 2^(-2*12) )   n = 12   d_n = -1-1i 
assign X[4'b1111] [13] = 144'h 000000000000200000000000012222221022;  // FFFFFFC00000080000 -0.0001220703112871 = 0.5 * ln( 1 + -1 * 2^(-13+1) + (-1^2+-1^2) * 2^(-2*13) )   n = 13   d_n = -1-1i 
assign X[4'b1111] [14] = 144'h 000000000000080000000000000488888884;  // FFFFFFE00000000000 -0.0000610351560984 = 0.5 * ln( 1 + -1 * 2^(-14+1) + (-1^2+-1^2) * 2^(-2*14) )   n = 14   d_n = -1-1i 
assign X[4'b1111] [15] = 144'h 000000000000020000000000000012222222;  // FFFFFFF00000000000 -0.0000305175781061 = 0.5 * ln( 1 + -1 * 2^(-15+1) + (-1^2+-1^2) * 2^(-2*15) )   n = 15   d_n = -1-1i 
assign X[4'b1111] [16] = 144'h 000000000000008000000000000000488888;  // FFFFFFF80000000000 -0.0000152587890601 = 0.5 * ln( 1 + -1 * 2^(-16+1) + (-1^2+-1^2) * 2^(-2*16) )   n = 16   d_n = -1-1i 
assign X[4'b1111] [17] = 144'h 000000000000002000000000000000012222;  // FFFFFFFC0000000000 -0.0000076293945310 = 0.5 * ln( 1 + -1 * 2^(-17+1) + (-1^2+-1^2) * 2^(-2*17) )   n = 17   d_n = -1-1i 
assign X[4'b1111] [18] = 144'h 000000000000000800000000000000000048;  // FFFFFFFE0000000000 -0.0000038146972656 = 0.5 * ln( 1 + -1 * 2^(-18+1) + (-1^2+-1^2) * 2^(-2*18) )   n = 18   d_n = -1-1i 
assign X[4'b1111] [19] = 144'h 000000000000000200000000000000000001;  // FFFFFFFF0000000000 -0.0000019073486328 = 0.5 * ln( 1 + -1 * 2^(-19+1) + (-1^2+-1^2) * 2^(-2*19) )   n = 19   d_n = -1-1i 
assign X[4'b1111] [20] = 144'h 000000000000000080000000000000000000;  // FFFFFFFF8000000000 -0.0000009536743164 = 0.5 * ln( 1 + -1 * 2^(-20+1) + (-1^2+-1^2) * 2^(-2*20) )   n = 20   d_n = -1-1i 
assign X[4'b1111] [21] = 144'h 000000000000000020000000000000000000;  // FFFFFFFFC000000000 -0.0000004768371582 = 0.5 * ln( 1 + -1 * 2^(-21+1) + (-1^2+-1^2) * 2^(-2*21) )   n = 21   d_n = -1-1i 
assign X[4'b1111] [22] = 144'h 000000000000000008000000000000000000;  // FFFFFFFFE000000000 -0.0000002384185791 = 0.5 * ln( 1 + -1 * 2^(-22+1) + (-1^2+-1^2) * 2^(-2*22) )   n = 22   d_n = -1-1i 
assign X[4'b1111] [23] = 144'h 000000000000000002000000000000000000;  // FFFFFFFFF000000000 -0.0000001192092896 = 0.5 * ln( 1 + -1 * 2^(-23+1) + (-1^2+-1^2) * 2^(-2*23) )   n = 23   d_n = -1-1i 
assign X[4'b1111] [24] = 144'h 000000000000000000800000000000000000;  // FFFFFFFFF800000000 -0.0000000596046448 = 0.5 * ln( 1 + -1 * 2^(-24+1) + (-1^2+-1^2) * 2^(-2*24) )   n = 24   d_n = -1-1i 
assign X[4'b1111] [25] = 144'h 000000000000000000200000000000000000;  // FFFFFFFFFC00000000 -0.0000000298023224 = 0.5 * ln( 1 + -1 * 2^(-25+1) + (-1^2+-1^2) * 2^(-2*25) )   n = 25   d_n = -1-1i 
assign X[4'b1111] [26] = 144'h 000000000000000000080000000000000000;  // FFFFFFFFFE00000000 -0.0000000149011612 = 0.5 * ln( 1 + -1 * 2^(-26+1) + (-1^2+-1^2) * 2^(-2*26) )   n = 26   d_n = -1-1i 
assign X[4'b1111] [27] = 144'h 000000000000000000020000000000000200;  // FFFFFFFFFF00000000 -0.0000000074505806 = 0.5 * ln( 1 + -1 * 2^(-27+1) + (-1^2+-1^2) * 2^(-2*27) )   n = 27   d_n = -1-1i 
assign X[4'b1111] [28] = 144'h 000000000000000000008000000000000020;  // FFFFFFFFFF80000000 -0.0000000037252903 = 0.5 * ln( 1 + -1 * 2^(-28+1) + (-1^2+-1^2) * 2^(-2*28) )   n = 28   d_n = -1-1i 
assign X[4'b1111] [29] = 144'h 000000000000000000002000000000000002;  // FFFFFFFFFFC0000000 -0.0000000018626452 = 0.5 * ln( 1 + -1 * 2^(-29+1) + (-1^2+-1^2) * 2^(-2*29) )   n = 29   d_n = -1-1i 
assign X[4'b1111] [30] = 144'h 000000000000000000000800000000000000;  // FFFFFFFFFFE0000000 -0.0000000009313226 = 0.5 * ln( 1 + -1 * 2^(-30+1) + (-1^2+-1^2) * 2^(-2*30) )   n = 30   d_n = -1-1i 
assign X[4'b1111] [31] = 144'h 000000000000000000000200000000000000;  // FFFFFFFFFFF0000000 -0.0000000004656613 = 0.5 * ln( 1 + -1 * 2^(-31+1) + (-1^2+-1^2) * 2^(-2*31) )   n = 31   d_n = -1-1i 
assign X[4'b1111] [32] = 144'h 000000000000000000000080000000000000;  // FFFFFFFFFFF8000000 -0.0000000002328306 = 0.5 * ln( 1 + -1 * 2^(-32+1) + (-1^2+-1^2) * 2^(-2*32) )   n = 32   d_n = -1-1i 
assign X[4'b1111] [33] = 144'h 000000000000000000000020000000000000;  // FFFFFFFFFFFC000000 -0.0000000001164153 = 0.5 * ln( 1 + -1 * 2^(-33+1) + (-1^2+-1^2) * 2^(-2*33) )   n = 33   d_n = -1-1i 
assign X[4'b1111] [34] = 144'h 000000000000000000000008000000000000;  // FFFFFFFFFFFE000000 -0.0000000000582077 = 0.5 * ln( 1 + -1 * 2^(-34+1) + (-1^2+-1^2) * 2^(-2*34) )   n = 34   d_n = -1-1i 
assign X[4'b1111] [35] = 144'h 000000000000000000000002000000000000;  // FFFFFFFFFFFF000000 -0.0000000000291038 = 0.5 * ln( 1 + -1 * 2^(-35+1) + (-1^2+-1^2) * 2^(-2*35) )   n = 35   d_n = -1-1i 
assign X[4'b1111] [36] = 144'h 000000000000000000000000800000000000;  // FFFFFFFFFFFF800000 -0.0000000000145519 = 0.5 * ln( 1 + -1 * 2^(-36+1) + (-1^2+-1^2) * 2^(-2*36) )   n = 36   d_n = -1-1i 
assign X[4'b1111] [37] = 144'h 000000000000000000000000200000000000;  // FFFFFFFFFFFFC00000 -0.0000000000072760 = 0.5 * ln( 1 + -1 * 2^(-37+1) + (-1^2+-1^2) * 2^(-2*37) )   n = 37   d_n = -1-1i 
assign X[4'b1111] [38] = 144'h 000000000000000000000000080000000000;  // FFFFFFFFFFFFE00000 -0.0000000000036380 = 0.5 * ln( 1 + -1 * 2^(-38+1) + (-1^2+-1^2) * 2^(-2*38) )   n = 38   d_n = -1-1i 
assign X[4'b1111] [39] = 144'h 000000000000000000000000020000000000;  // FFFFFFFFFFFFF00000 -0.0000000000018190 = 0.5 * ln( 1 + -1 * 2^(-39+1) + (-1^2+-1^2) * 2^(-2*39) )   n = 39   d_n = -1-1i 
assign X[4'b1111] [40] = 144'h 000000000000000000000000008000000000;  // FFFFFFFFFFFFF80000 -0.0000000000009095 = 0.5 * ln( 1 + -1 * 2^(-40+1) + (-1^2+-1^2) * 2^(-2*40) )   n = 40   d_n = -1-1i 
assign X[4'b1111] [41] = 144'h 000000000000000000000000002000000000;  // FFFFFFFFFFFFF80000 -0.0000000000004547 = 0.5 * ln( 1 + -1 * 2^(-41+1) + (-1^2+-1^2) * 2^(-2*41) )   n = 41   d_n = -1-1i 
assign X[4'b1111] [42] = 144'h 000000000000000000000000000800000000;  // 1000000000000000000 -0.0000000000002274 = 0.5 * ln( 1 + -1 * 2^(-42+1) + (-1^2+-1^2) * 2^(-2*42) )   n = 42   d_n = -1-1i 
assign X[4'b1111] [43] = 144'h 000000000000000000000000000200000000;  // 1000000000000000000 -0.0000000000001137 = 0.5 * ln( 1 + -1 * 2^(-43+1) + (-1^2+-1^2) * 2^(-2*43) )   n = 43   d_n = -1-1i 
assign X[4'b1111] [44] = 144'h 000000000000000000000000000080000000;  // 1000000000000000000 -0.0000000000000568 = 0.5 * ln( 1 + -1 * 2^(-44+1) + (-1^2+-1^2) * 2^(-2*44) )   n = 44   d_n = -1-1i 
assign X[4'b1111] [45] = 144'h 000000000000000000000000000020000000;  // 1000000000000000000 -0.0000000000000284 = 0.5 * ln( 1 + -1 * 2^(-45+1) + (-1^2+-1^2) * 2^(-2*45) )   n = 45   d_n = -1-1i 
assign X[4'b1111] [46] = 144'h 000000000000000000000000000008000000;  // 1000000000000000000 -0.0000000000000142 = 0.5 * ln( 1 + -1 * 2^(-46+1) + (-1^2+-1^2) * 2^(-2*46) )   n = 46   d_n = -1-1i 
assign X[4'b1111] [47] = 144'h 000000000000000000000000000002000000;  // 1000000000000000000 -0.0000000000000071 = 0.5 * ln( 1 + -1 * 2^(-47+1) + (-1^2+-1^2) * 2^(-2*47) )   n = 47   d_n = -1-1i 
assign X[4'b1111] [48] = 144'h 000000000000000000000000000000800000;  // 1000000000000000000 -0.0000000000000036 = 0.5 * ln( 1 + -1 * 2^(-48+1) + (-1^2+-1^2) * 2^(-2*48) )   n = 48   d_n = -1-1i 
assign X[4'b1111] [49] = 144'h 000000000000000000000000000000200000;  // 1000000000000000000 -0.0000000000000018 = 0.5 * ln( 1 + -1 * 2^(-49+1) + (-1^2+-1^2) * 2^(-2*49) )   n = 49   d_n = -1-1i 
assign X[4'b1111] [50] = 144'h 000000000000000000000000000000080000;  // 1000000000000000000 -0.0000000000000009 = 0.5 * ln( 1 + -1 * 2^(-50+1) + (-1^2+-1^2) * 2^(-2*50) )   n = 50   d_n = -1-1i 
assign X[4'b1111] [51] = 144'h 000000000000000000000000000000020000;  // 1000000000000000000 -0.0000000000000004 = 0.5 * ln( 1 + -1 * 2^(-51+1) + (-1^2+-1^2) * 2^(-2*51) )   n = 51   d_n = -1-1i 
assign X[4'b1111] [52] = 144'h 000000000000000000000000000000008000;  // 1000000000000000000 -0.0000000000000002 = 0.5 * ln( 1 + -1 * 2^(-52+1) + (-1^2+-1^2) * 2^(-2*52) )   n = 52   d_n = -1-1i 
assign X[4'b1111] [53] = 144'h 000000000000000000000000000000002000;  // 1000000000000000000 -0.0000000000000001 = 0.5 * ln( 1 + -1 * 2^(-53+1) + (-1^2+-1^2) * 2^(-2*53) )   n = 53   d_n = -1-1i 
assign X[4'b1111] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-54+1) + (-1^2+-1^2) * 2^(-2*54) )   n = 54   d_n = -1-1i 
assign X[4'b1111] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-55+1) + (-1^2+-1^2) * 2^(-2*55) )   n = 55   d_n = -1-1i 
assign X[4'b1111] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-56+1) + (-1^2+-1^2) * 2^(-2*56) )   n = 56   d_n = -1-1i 
assign X[4'b1111] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-57+1) + (-1^2+-1^2) * 2^(-2*57) )   n = 57   d_n = -1-1i 
assign X[4'b1111] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-58+1) + (-1^2+-1^2) * 2^(-2*58) )   n = 58   d_n = -1-1i 
assign X[4'b1111] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-59+1) + (-1^2+-1^2) * 2^(-2*59) )   n = 59   d_n = -1-1i 
assign X[4'b1111] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-60+1) + (-1^2+-1^2) * 2^(-2*60) )   n = 60   d_n = -1-1i 
assign X[4'b1111] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-61+1) + (-1^2+-1^2) * 2^(-2*61) )   n = 61   d_n = -1-1i 
assign X[4'b1111] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-62+1) + (-1^2+-1^2) * 2^(-2*62) )   n = 62   d_n = -1-1i 
assign X[4'b1111] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-63+1) + (-1^2+-1^2) * 2^(-2*63) )   n = 63   d_n = -1-1i 
assign X[4'b1111] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 = 0.5 * ln( 1 + -1 * 2^(-64+1) + (-1^2+-1^2) * 2^(-2*64) )   n = 64   d_n = -1-1i 
assign Y[4'b0000] [01] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = 0 
assign Y[4'b0000] [02] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = 0 
assign Y[4'b0000] [03] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = 0 
assign Y[4'b0000] [04] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = 0 
assign Y[4'b0000] [05] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = 0 
assign Y[4'b0000] [06] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = 0 
assign Y[4'b0000] [07] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = 0 
assign Y[4'b0000] [08] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = 0 
assign Y[4'b0000] [09] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = 0 
assign Y[4'b0000] [10] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = 0 
assign Y[4'b0000] [11] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = 0 
assign Y[4'b0000] [12] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = 0 
assign Y[4'b0000] [13] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = 0 
assign Y[4'b0000] [14] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = 0 
assign Y[4'b0000] [15] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = 0 
assign Y[4'b0000] [16] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = 0 
assign Y[4'b0000] [17] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = 0 
assign Y[4'b0000] [18] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = 0 
assign Y[4'b0000] [19] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = 0 
assign Y[4'b0000] [20] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = 0 
assign Y[4'b0000] [21] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = 0 
assign Y[4'b0000] [22] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = 0 
assign Y[4'b0000] [23] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = 0 
assign Y[4'b0000] [24] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = 0 
assign Y[4'b0000] [25] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = 0 
assign Y[4'b0000] [26] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = 0 
assign Y[4'b0000] [27] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = 0 
assign Y[4'b0000] [28] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = 0 
assign Y[4'b0000] [29] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = 0 
assign Y[4'b0000] [30] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = 0 
assign Y[4'b0000] [31] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = 0 
assign Y[4'b0000] [32] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = 0 
assign Y[4'b0000] [33] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = 0 
assign Y[4'b0000] [34] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = 0 
assign Y[4'b0000] [35] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = 0 
assign Y[4'b0000] [36] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = 0 
assign Y[4'b0000] [37] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = 0 
assign Y[4'b0000] [38] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = 0 
assign Y[4'b0000] [39] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = 0 
assign Y[4'b0000] [40] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = 0 
assign Y[4'b0000] [41] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = 0 
assign Y[4'b0000] [42] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = 0 
assign Y[4'b0000] [43] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = 0 
assign Y[4'b0000] [44] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = 0 
assign Y[4'b0000] [45] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = 0 
assign Y[4'b0000] [46] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = 0 
assign Y[4'b0000] [47] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = 0 
assign Y[4'b0000] [48] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = 0 
assign Y[4'b0000] [49] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = 0 
assign Y[4'b0000] [50] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = 0 
assign Y[4'b0000] [51] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = 0 
assign Y[4'b0000] [52] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = 0 
assign Y[4'b0000] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = 0 
assign Y[4'b0000] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = 0 
assign Y[4'b0000] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = 0 
assign Y[4'b0000] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = 0 
assign Y[4'b0000] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = 0 
assign Y[4'b0000] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = 0 
assign Y[4'b0000] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = 0 
assign Y[4'b0000] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = 0 
assign Y[4'b0000] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = 0 
assign Y[4'b0000] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = 0 
assign Y[4'b0000] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = 0 
assign Y[4'b0000] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = 0 
assign Y[4'b0001] [01] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^1 ) )   n =  1   d_n = 1 
assign Y[4'b0001] [02] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^2 ) )   n =  2   d_n = 1 
assign Y[4'b0001] [03] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^3 ) )   n =  3   d_n = 1 
assign Y[4'b0001] [04] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^4 ) )   n =  4   d_n = 1 
assign Y[4'b0001] [05] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^5 ) )   n =  5   d_n = 1 
assign Y[4'b0001] [06] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^6 ) )   n =  6   d_n = 1 
assign Y[4'b0001] [07] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^7 ) )   n =  7   d_n = 1 
assign Y[4'b0001] [08] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^8 ) )   n =  8   d_n = 1 
assign Y[4'b0001] [09] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^9 ) )   n =  9   d_n = 1 
assign Y[4'b0001] [10] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^10 ) )   n = 10   d_n = 1 
assign Y[4'b0001] [11] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^11 ) )   n = 11   d_n = 1 
assign Y[4'b0001] [12] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^12 ) )   n = 12   d_n = 1 
assign Y[4'b0001] [13] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^13 ) )   n = 13   d_n = 1 
assign Y[4'b0001] [14] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^14 ) )   n = 14   d_n = 1 
assign Y[4'b0001] [15] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^15 ) )   n = 15   d_n = 1 
assign Y[4'b0001] [16] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^16 ) )   n = 16   d_n = 1 
assign Y[4'b0001] [17] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^17 ) )   n = 17   d_n = 1 
assign Y[4'b0001] [18] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^18 ) )   n = 18   d_n = 1 
assign Y[4'b0001] [19] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^19 ) )   n = 19   d_n = 1 
assign Y[4'b0001] [20] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^20 ) )   n = 20   d_n = 1 
assign Y[4'b0001] [21] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^21 ) )   n = 21   d_n = 1 
assign Y[4'b0001] [22] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^22 ) )   n = 22   d_n = 1 
assign Y[4'b0001] [23] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^23 ) )   n = 23   d_n = 1 
assign Y[4'b0001] [24] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^24 ) )   n = 24   d_n = 1 
assign Y[4'b0001] [25] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^25 ) )   n = 25   d_n = 1 
assign Y[4'b0001] [26] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^26 ) )   n = 26   d_n = 1 
assign Y[4'b0001] [27] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^27 ) )   n = 27   d_n = 1 
assign Y[4'b0001] [28] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^28 ) )   n = 28   d_n = 1 
assign Y[4'b0001] [29] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^29 ) )   n = 29   d_n = 1 
assign Y[4'b0001] [30] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^30 ) )   n = 30   d_n = 1 
assign Y[4'b0001] [31] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^31 ) )   n = 31   d_n = 1 
assign Y[4'b0001] [32] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^32 ) )   n = 32   d_n = 1 
assign Y[4'b0001] [33] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^33 ) )   n = 33   d_n = 1 
assign Y[4'b0001] [34] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^34 ) )   n = 34   d_n = 1 
assign Y[4'b0001] [35] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^35 ) )   n = 35   d_n = 1 
assign Y[4'b0001] [36] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^36 ) )   n = 36   d_n = 1 
assign Y[4'b0001] [37] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^37 ) )   n = 37   d_n = 1 
assign Y[4'b0001] [38] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^38 ) )   n = 38   d_n = 1 
assign Y[4'b0001] [39] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^39 ) )   n = 39   d_n = 1 
assign Y[4'b0001] [40] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^40 ) )   n = 40   d_n = 1 
assign Y[4'b0001] [41] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^41 ) )   n = 41   d_n = 1 
assign Y[4'b0001] [42] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^42 ) )   n = 42   d_n = 1 
assign Y[4'b0001] [43] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^43 ) )   n = 43   d_n = 1 
assign Y[4'b0001] [44] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^44 ) )   n = 44   d_n = 1 
assign Y[4'b0001] [45] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^45 ) )   n = 45   d_n = 1 
assign Y[4'b0001] [46] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^46 ) )   n = 46   d_n = 1 
assign Y[4'b0001] [47] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^47 ) )   n = 47   d_n = 1 
assign Y[4'b0001] [48] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^48 ) )   n = 48   d_n = 1 
assign Y[4'b0001] [49] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^49 ) )   n = 49   d_n = 1 
assign Y[4'b0001] [50] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^50 ) )   n = 50   d_n = 1 
assign Y[4'b0001] [51] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^51 ) )   n = 51   d_n = 1 
assign Y[4'b0001] [52] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^52 ) )   n = 52   d_n = 1 
assign Y[4'b0001] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^53 ) )   n = 53   d_n = 1 
assign Y[4'b0001] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^54 ) )   n = 54   d_n = 1 
assign Y[4'b0001] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^55 ) )   n = 55   d_n = 1 
assign Y[4'b0001] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^56 ) )   n = 56   d_n = 1 
assign Y[4'b0001] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^57 ) )   n = 57   d_n = 1 
assign Y[4'b0001] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^58 ) )   n = 58   d_n = 1 
assign Y[4'b0001] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^59 ) )   n = 59   d_n = 1 
assign Y[4'b0001] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^60 ) )   n = 60   d_n = 1 
assign Y[4'b0001] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^61 ) )   n = 61   d_n = 1 
assign Y[4'b0001] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^62 ) )   n = 62   d_n = 1 
assign Y[4'b0001] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^63 ) )   n = 63   d_n = 1 
assign Y[4'b0001] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^64 ) )   n = 64   d_n = 1 
assign Y[4'b0010] [01] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = -0 
assign Y[4'b0010] [02] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = -0 
assign Y[4'b0010] [03] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = -0 
assign Y[4'b0010] [04] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = -0 
assign Y[4'b0010] [05] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = -0 
assign Y[4'b0010] [06] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = -0 
assign Y[4'b0010] [07] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = -0 
assign Y[4'b0010] [08] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = -0 
assign Y[4'b0010] [09] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = -0 
assign Y[4'b0010] [10] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = -0 
assign Y[4'b0010] [11] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = -0 
assign Y[4'b0010] [12] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = -0 
assign Y[4'b0010] [13] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = -0 
assign Y[4'b0010] [14] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = -0 
assign Y[4'b0010] [15] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = -0 
assign Y[4'b0010] [16] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = -0 
assign Y[4'b0010] [17] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = -0 
assign Y[4'b0010] [18] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = -0 
assign Y[4'b0010] [19] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = -0 
assign Y[4'b0010] [20] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = -0 
assign Y[4'b0010] [21] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = -0 
assign Y[4'b0010] [22] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = -0 
assign Y[4'b0010] [23] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = -0 
assign Y[4'b0010] [24] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = -0 
assign Y[4'b0010] [25] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = -0 
assign Y[4'b0010] [26] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = -0 
assign Y[4'b0010] [27] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = -0 
assign Y[4'b0010] [28] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = -0 
assign Y[4'b0010] [29] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = -0 
assign Y[4'b0010] [30] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = -0 
assign Y[4'b0010] [31] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = -0 
assign Y[4'b0010] [32] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = -0 
assign Y[4'b0010] [33] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = -0 
assign Y[4'b0010] [34] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = -0 
assign Y[4'b0010] [35] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = -0 
assign Y[4'b0010] [36] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = -0 
assign Y[4'b0010] [37] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = -0 
assign Y[4'b0010] [38] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = -0 
assign Y[4'b0010] [39] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = -0 
assign Y[4'b0010] [40] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = -0 
assign Y[4'b0010] [41] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = -0 
assign Y[4'b0010] [42] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = -0 
assign Y[4'b0010] [43] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = -0 
assign Y[4'b0010] [44] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = -0 
assign Y[4'b0010] [45] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = -0 
assign Y[4'b0010] [46] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = -0 
assign Y[4'b0010] [47] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = -0 
assign Y[4'b0010] [48] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = -0 
assign Y[4'b0010] [49] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = -0 
assign Y[4'b0010] [50] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = -0 
assign Y[4'b0010] [51] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = -0 
assign Y[4'b0010] [52] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = -0 
assign Y[4'b0010] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = -0 
assign Y[4'b0010] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = -0 
assign Y[4'b0010] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = -0 
assign Y[4'b0010] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = -0 
assign Y[4'b0010] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = -0 
assign Y[4'b0010] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = -0 
assign Y[4'b0010] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = -0 
assign Y[4'b0010] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = -0 
assign Y[4'b0010] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = -0 
assign Y[4'b0010] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = -0 
assign Y[4'b0010] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = -0 
assign Y[4'b0010] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = -0 
assign Y[4'b0011] [01] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^1 ) )   n =  1   d_n = -1 
assign Y[4'b0011] [02] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^2 ) )   n =  2   d_n = -1 
assign Y[4'b0011] [03] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^3 ) )   n =  3   d_n = -1 
assign Y[4'b0011] [04] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^4 ) )   n =  4   d_n = -1 
assign Y[4'b0011] [05] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^5 ) )   n =  5   d_n = -1 
assign Y[4'b0011] [06] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^6 ) )   n =  6   d_n = -1 
assign Y[4'b0011] [07] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^7 ) )   n =  7   d_n = -1 
assign Y[4'b0011] [08] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^8 ) )   n =  8   d_n = -1 
assign Y[4'b0011] [09] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^9 ) )   n =  9   d_n = -1 
assign Y[4'b0011] [10] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^10 ) )   n = 10   d_n = -1 
assign Y[4'b0011] [11] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^11 ) )   n = 11   d_n = -1 
assign Y[4'b0011] [12] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^12 ) )   n = 12   d_n = -1 
assign Y[4'b0011] [13] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^13 ) )   n = 13   d_n = -1 
assign Y[4'b0011] [14] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^14 ) )   n = 14   d_n = -1 
assign Y[4'b0011] [15] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^15 ) )   n = 15   d_n = -1 
assign Y[4'b0011] [16] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^16 ) )   n = 16   d_n = -1 
assign Y[4'b0011] [17] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^17 ) )   n = 17   d_n = -1 
assign Y[4'b0011] [18] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^18 ) )   n = 18   d_n = -1 
assign Y[4'b0011] [19] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^19 ) )   n = 19   d_n = -1 
assign Y[4'b0011] [20] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^20 ) )   n = 20   d_n = -1 
assign Y[4'b0011] [21] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^21 ) )   n = 21   d_n = -1 
assign Y[4'b0011] [22] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^22 ) )   n = 22   d_n = -1 
assign Y[4'b0011] [23] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^23 ) )   n = 23   d_n = -1 
assign Y[4'b0011] [24] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^24 ) )   n = 24   d_n = -1 
assign Y[4'b0011] [25] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^25 ) )   n = 25   d_n = -1 
assign Y[4'b0011] [26] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^26 ) )   n = 26   d_n = -1 
assign Y[4'b0011] [27] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^27 ) )   n = 27   d_n = -1 
assign Y[4'b0011] [28] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^28 ) )   n = 28   d_n = -1 
assign Y[4'b0011] [29] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^29 ) )   n = 29   d_n = -1 
assign Y[4'b0011] [30] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^30 ) )   n = 30   d_n = -1 
assign Y[4'b0011] [31] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^31 ) )   n = 31   d_n = -1 
assign Y[4'b0011] [32] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^32 ) )   n = 32   d_n = -1 
assign Y[4'b0011] [33] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^33 ) )   n = 33   d_n = -1 
assign Y[4'b0011] [34] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^34 ) )   n = 34   d_n = -1 
assign Y[4'b0011] [35] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^35 ) )   n = 35   d_n = -1 
assign Y[4'b0011] [36] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^36 ) )   n = 36   d_n = -1 
assign Y[4'b0011] [37] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^37 ) )   n = 37   d_n = -1 
assign Y[4'b0011] [38] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^38 ) )   n = 38   d_n = -1 
assign Y[4'b0011] [39] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^39 ) )   n = 39   d_n = -1 
assign Y[4'b0011] [40] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^40 ) )   n = 40   d_n = -1 
assign Y[4'b0011] [41] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^41 ) )   n = 41   d_n = -1 
assign Y[4'b0011] [42] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^42 ) )   n = 42   d_n = -1 
assign Y[4'b0011] [43] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^43 ) )   n = 43   d_n = -1 
assign Y[4'b0011] [44] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^44 ) )   n = 44   d_n = -1 
assign Y[4'b0011] [45] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^45 ) )   n = 45   d_n = -1 
assign Y[4'b0011] [46] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^46 ) )   n = 46   d_n = -1 
assign Y[4'b0011] [47] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^47 ) )   n = 47   d_n = -1 
assign Y[4'b0011] [48] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^48 ) )   n = 48   d_n = -1 
assign Y[4'b0011] [49] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^49 ) )   n = 49   d_n = -1 
assign Y[4'b0011] [50] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^50 ) )   n = 50   d_n = -1 
assign Y[4'b0011] [51] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^51 ) )   n = 51   d_n = -1 
assign Y[4'b0011] [52] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^52 ) )   n = 52   d_n = -1 
assign Y[4'b0011] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^53 ) )   n = 53   d_n = -1 
assign Y[4'b0011] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^54 ) )   n = 54   d_n = -1 
assign Y[4'b0011] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^55 ) )   n = 55   d_n = -1 
assign Y[4'b0011] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^56 ) )   n = 56   d_n = -1 
assign Y[4'b0011] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^57 ) )   n = 57   d_n = -1 
assign Y[4'b0011] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^58 ) )   n = 58   d_n = -1 
assign Y[4'b0011] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^59 ) )   n = 59   d_n = -1 
assign Y[4'b0011] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^60 ) )   n = 60   d_n = -1 
assign Y[4'b0011] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^61 ) )   n = 61   d_n = -1 
assign Y[4'b0011] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^62 ) )   n = 62   d_n = -1 
assign Y[4'b0011] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^63 ) )   n = 63   d_n = -1 
assign Y[4'b0011] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^64 ) )   n = 64   d_n = -1 
assign Y[4'b0100] [01] = 144'h 000000102088812108012220108088440800;  // 0003B58CE0AC3769E0 +0.4636476090008061 =  1 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = 0+1i 
assign Y[4'b0100] [02] = 144'h 000000040088208088008112204001082000;  // 0001F5B75F92C80DD0 +0.2449786631268641 =  1 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = 0+1i 
assign Y[4'b0100] [03] = 144'h 000000010002220821110888880480208200;  // 0000FEADD4D5617B70 +0.1243549945467614 =  1 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = 0+1i 
assign Y[4'b0100] [04] = 144'h 000000004000088882020821221000808440;  // 00007FD56EDCB3F7A8 +0.0624188099959574 =  1 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = 0+1i 
assign Y[4'b0100] [05] = 144'h 000000001000002222208082111202201040;  // 00003FFAAB7752EC4A +0.0312398334302683 =  1 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = 0+1i 
assign Y[4'b0100] [06] = 144'h 000000000400000088888820202082044422;  // 00001FFF555BBB729B +0.0156237286204768 =  1 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = 0+1i 
assign Y[4'b0100] [07] = 144'h 000000000100000002222222080808211120;  // 00000FFFEAAADDDD4B +0.0078123410601011 =  1 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = 0+1i 
assign Y[4'b0100] [08] = 144'h 000000000040000000088888888202020208;  // 000007FFFD5556EEED +0.0039062301319670 =  1 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = 0+1i 
assign Y[4'b0100] [09] = 144'h 000000000010000000002222222220808080;  // 000003FFFFAAAAB777 +0.0019531225164788 =  1 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = 0+1i 
assign Y[4'b0100] [10] = 144'h 000000000004000000000088888888882020;  // 000001FFFFF55555BB +0.0009765621895593 =  1 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = 0+1i 
assign Y[4'b0100] [11] = 144'h 000000000001000000000002222222222208;  // 000000FFFFFEAAAAAD +0.0004882812111949 =  1 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = 0+1i 
assign Y[4'b0100] [12] = 144'h 000000000000400000000000088888888888;  // 0000007FFFFFD55555 +0.0002441406201494 =  1 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = 0+1i 
assign Y[4'b0100] [13] = 144'h 000000000000100000000000008444444444;  // 0000003FFFFFFAAAAA +0.0001220703118937 =  1 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = 0+1i 
assign Y[4'b0100] [14] = 144'h 000000000000040000000000000211111111;  // 0000001FFFFFFF5555 +0.0000610351561742 =  1 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = 0+1i 
assign Y[4'b0100] [15] = 144'h 000000000000010000000000000008444444;  // 0000000FFFFFFFEAAA +0.0000305175781155 =  1 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = 0+1i 
assign Y[4'b0100] [16] = 144'h 000000000000004000000000000000211111;  // 00000007FFFFFFFD55 +0.0000152587890613 =  1 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = 0+1i 
assign Y[4'b0100] [17] = 144'h 000000000000001000000000000000008444;  // 00000003FFFFFFFFAA +0.0000076293945311 =  1 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = 0+1i 
assign Y[4'b0100] [18] = 144'h 000000000000000400000000000000000211;  // 00000001FFFFFFFFF5 +0.0000038146972656 =  1 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = 0+1i 
assign Y[4'b0100] [19] = 144'h 000000000000000100000000000000000008;  // 00000000FFFFFFFFFE +0.0000019073486328 =  1 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = 0+1i 
assign Y[4'b0100] [20] = 144'h 000000000000000040000000000000000000;  // 000000007FFFFFFFFF +0.0000009536743164 =  1 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = 0+1i 
assign Y[4'b0100] [21] = 144'h 000000000000000010000000000000000000;  // 000000003FFFFFFFFF +0.0000004768371582 =  1 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = 0+1i 
assign Y[4'b0100] [22] = 144'h 000000000000000004000000000000000000;  // 000000001FFFFFFFFF +0.0000002384185791 =  1 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = 0+1i 
assign Y[4'b0100] [23] = 144'h 000000000000000001000000000000000000;  // 000000000FFFFFFFFF +0.0000001192092896 =  1 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = 0+1i 
assign Y[4'b0100] [24] = 144'h 000000000000000000400000000000000000;  // 0000000007FFFFFFFF +0.0000000596046448 =  1 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = 0+1i 
assign Y[4'b0100] [25] = 144'h 000000000000000000100000000000000000;  // 0000000003FFFFFFFF +0.0000000298023224 =  1 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = 0+1i 
assign Y[4'b0100] [26] = 144'h 000000000000000000040000000000000000;  // 0000000001FFFFFFFF +0.0000000149011612 =  1 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = 0+1i 
assign Y[4'b0100] [27] = 144'h 000000000000000000010000000000000000;  // 000000000100000000 +0.0000000074505806 =  1 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = 0+1i 
assign Y[4'b0100] [28] = 144'h 000000000000000000004000000000000000;  // 000000000080000000 +0.0000000037252903 =  1 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = 0+1i 
assign Y[4'b0100] [29] = 144'h 000000000000000000001000000000000000;  // 000000000040000000 +0.0000000018626451 =  1 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = 0+1i 
assign Y[4'b0100] [30] = 144'h 000000000000000000000400000000000000;  // 000000000020000000 +0.0000000009313226 =  1 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = 0+1i 
assign Y[4'b0100] [31] = 144'h 000000000000000000000100000000000000;  // 000000000010000000 +0.0000000004656613 =  1 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = 0+1i 
assign Y[4'b0100] [32] = 144'h 000000000000000000000040000000000000;  // 000000000008000000 +0.0000000002328306 =  1 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = 0+1i 
assign Y[4'b0100] [33] = 144'h 000000000000000000000010000000000000;  // 000000000004000000 +0.0000000001164153 =  1 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = 0+1i 
assign Y[4'b0100] [34] = 144'h 000000000000000000000004000000000000;  // 000000000002000000 +0.0000000000582077 =  1 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = 0+1i 
assign Y[4'b0100] [35] = 144'h 000000000000000000000001000000000000;  // 000000000001000000 +0.0000000000291038 =  1 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = 0+1i 
assign Y[4'b0100] [36] = 144'h 000000000000000000000000400000000000;  // 000000000000800000 +0.0000000000145519 =  1 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = 0+1i 
assign Y[4'b0100] [37] = 144'h 000000000000000000000000100000000000;  // 000000000000400000 +0.0000000000072760 =  1 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = 0+1i 
assign Y[4'b0100] [38] = 144'h 000000000000000000000000040000000000;  // 000000000000200000 +0.0000000000036380 =  1 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = 0+1i 
assign Y[4'b0100] [39] = 144'h 000000000000000000000000010000000000;  // 000000000000100000 +0.0000000000018190 =  1 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = 0+1i 
assign Y[4'b0100] [40] = 144'h 000000000000000000000000004000000000;  // 000000000000080000 +0.0000000000009095 =  1 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = 0+1i 
assign Y[4'b0100] [41] = 144'h 000000000000000000000000001000000000;  // 000000000000040000 +0.0000000000004547 =  1 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = 0+1i 
assign Y[4'b0100] [42] = 144'h 000000000000000000000000000400000000;  // 000000000000020000 +0.0000000000002274 =  1 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = 0+1i 
assign Y[4'b0100] [43] = 144'h 000000000000000000000000000100000000;  // 000000000000010000 +0.0000000000001137 =  1 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = 0+1i 
assign Y[4'b0100] [44] = 144'h 000000000000000000000000000040000000;  // 000000000000008000 +0.0000000000000568 =  1 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = 0+1i 
assign Y[4'b0100] [45] = 144'h 000000000000000000000000000010000000;  // 000000000000004000 +0.0000000000000284 =  1 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = 0+1i 
assign Y[4'b0100] [46] = 144'h 000000000000000000000000000004000000;  // 000000000000002000 +0.0000000000000142 =  1 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = 0+1i 
assign Y[4'b0100] [47] = 144'h 000000000000000000000000000001000000;  // 000000000000001000 +0.0000000000000071 =  1 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = 0+1i 
assign Y[4'b0100] [48] = 144'h 000000000000000000000000000000400000;  // 000000000000000800 +0.0000000000000036 =  1 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = 0+1i 
assign Y[4'b0100] [49] = 144'h 000000000000000000000000000000100000;  // 000000000000000400 +0.0000000000000018 =  1 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = 0+1i 
assign Y[4'b0100] [50] = 144'h 000000000000000000000000000000040000;  // 000000000000000200 +0.0000000000000009 =  1 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = 0+1i 
assign Y[4'b0100] [51] = 144'h 000000000000000000000000000000010000;  // 000000000000000100 +0.0000000000000004 =  1 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = 0+1i 
assign Y[4'b0100] [52] = 144'h 000000000000000000000000000000004000;  // 000000000000000080 +0.0000000000000002 =  1 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = 0+1i 
assign Y[4'b0100] [53] = 144'h 000000000000000000000000000000001000;  // 000000000000000040 +0.0000000000000001 =  1 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = 0+1i 
assign Y[4'b0100] [54] = 144'h 000000000000000000000000000000000400;  // 000000000000000020 +0.0000000000000001 =  1 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = 0+1i 
assign Y[4'b0100] [55] = 144'h 000000000000000000000000000000000100;  // 000000000000000010 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = 0+1i 
assign Y[4'b0100] [56] = 144'h 000000000000000000000000000000000040;  // 000000000000000008 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = 0+1i 
assign Y[4'b0100] [57] = 144'h 000000000000000000000000000000000010;  // 000000000000000004 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = 0+1i 
assign Y[4'b0100] [58] = 144'h 000000000000000000000000000000000004;  // 000000000000000002 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = 0+1i 
assign Y[4'b0100] [59] = 144'h 000000000000000000000000000000000001;  // 000000000000000001 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = 0+1i 
assign Y[4'b0100] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = 0+1i 
assign Y[4'b0100] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = 0+1i 
assign Y[4'b0100] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = 0+1i 
assign Y[4'b0100] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = 0+1i 
assign Y[4'b0100] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = 0+1i 
assign Y[4'b0101] [01] = 144'h 000000044112020402104811211008200400;  // 000292F1F464D3DC20 +0.3217505543966422 =  1 * atan( 1 / (  1 + 2^1 ) )   n =  1   d_n = 1+1i 
assign Y[4'b0101] [02] = 144'h 000000048110101004008100820448012200;  // 000194441F8F7260B0 +0.1973955598498807 =  1 * atan( 1 / (  1 + 2^2 ) )   n =  2   d_n = 1+1i 
assign Y[4'b0101] [03] = 144'h 000000010804440010012100010044048000;  // 0000E2A040D010A180 +0.1106572211738956 =  1 * atan( 1 / (  1 + 2^3 ) )   n =  3   d_n = 1+1i 
assign Y[4'b0101] [04] = 144'h 000000004080111100810040042008202100;  // 00007854F9081BDBD4 +0.0587558227157227 =  1 * atan( 1 / (  1 + 2^4 ) )   n =  4   d_n = 1+1i 
assign Y[4'b0101] [05] = 144'h 000000001008004444408401000800208840;  // 00003E0AA7A0FDFB68 +0.0302937599187751 =  1 * atan( 1 / (  1 + 2^5 ) )   n =  5   d_n = 1+1i 
assign Y[4'b0101] [06] = 144'h 000000000400800111111020481004088080;  // 00001F81553C641D79 +0.0153834017805952 =  1 * atan( 1 / (  1 + 2^6 ) )   n =  6   d_n = 1+1i 
assign Y[4'b0101] [07] = 144'h 000000000100080004444444080040100088;  // 00000FE02AA9E083F6 +0.0077517827122069 =  1 * atan( 1 / (  1 + 2^7 ) )   n =  7   d_n = 1+1i 
assign Y[4'b0101] [08] = 144'h 000000000040008000111111110200848100;  // 000007F805554EF990 +0.0038910309466445 =  1 * atan( 1 / (  1 + 2^8 ) )   n =  8   d_n = 1+1i 
assign Y[4'b0101] [09] = 144'h 000000000010000800004444444440808404;  // 000003FE00AAAA77A2 +0.0019493152697654 =  1 * atan( 1 / (  1 + 2^9 ) )   n =  9   d_n = 1+1i 
assign Y[4'b0101] [10] = 144'h 000000000004000080000111111111102020;  // 000001FF80155553BC +0.0009756094465646 =  1 * atan( 1 / (  1 + 2^10 ) )   n = 10   d_n = 1+1i 
assign Y[4'b0101] [11] = 144'h 000000000001000008000004444444444408;  // 000000FFE002AAAA9D +0.0004880429090311 =  1 * atan( 1 / (  1 + 2^11 ) )   n = 11   d_n = 1+1i 
assign Y[4'b0101] [12] = 144'h 000000000000400000800000111111111111;  // 0000007FF800555554 +0.0002440810300565 =  1 * atan( 1 / (  1 + 2^12 ) )   n = 12   d_n = 1+1i 
assign Y[4'b0101] [13] = 144'h 000000000000100000080000004444444444;  // 0000003FFE000AAAAA +0.0001220554125515 =  1 * atan( 1 / (  1 + 2^13 ) )   n = 13   d_n = 1+1i 
assign Y[4'b0101] [14] = 144'h 000000000000040000008000000111111111;  // 0000001FFF80015555 +0.0000610314311113 =  1 * atan( 1 / (  1 + 2^14 ) )   n = 14   d_n = 1+1i 
assign Y[4'b0101] [15] = 144'h 000000000000010000000800000004444444;  // 0000000FFFE0002AAA +0.0000305166468214 =  1 * atan( 1 / (  1 + 2^15 ) )   n = 15   d_n = 1+1i 
assign Y[4'b0101] [16] = 144'h 000000000000004000000080000000111111;  // 00000007FFF8000555 +0.0000152585562342 =  1 * atan( 1 / (  1 + 2^16 ) )   n = 16   d_n = 1+1i 
assign Y[4'b0101] [17] = 144'h 000000000000001000000008000000004444;  // 00000003FFFE0000AA +0.0000076293363239 =  1 * atan( 1 / (  1 + 2^17 ) )   n = 17   d_n = 1+1i 
assign Y[4'b0101] [18] = 144'h 000000000000000400000000800000000111;  // 00000001FFFF800015 +0.0000038146827137 =  1 * atan( 1 / (  1 + 2^18 ) )   n = 18   d_n = 1+1i 
assign Y[4'b0101] [19] = 144'h 000000000000000100000000080000000004;  // 00000000FFFFE00002 +0.0000019073449948 =  1 * atan( 1 / (  1 + 2^19 ) )   n = 19   d_n = 1+1i 
assign Y[4'b0101] [20] = 144'h 000000000000000040000000008000000000;  // 000000007FFFF80000 +0.0000009536734069 =  1 * atan( 1 / (  1 + 2^20 ) )   n = 20   d_n = 1+1i 
assign Y[4'b0101] [21] = 144'h 000000000000000010000000000800000000;  // 000000003FFFFE0000 +0.0000004768369308 =  1 * atan( 1 / (  1 + 2^21 ) )   n = 21   d_n = 1+1i 
assign Y[4'b0101] [22] = 144'h 000000000000000004000000000080000000;  // 000000001FFFFF8000 +0.0000002384185223 =  1 * atan( 1 / (  1 + 2^22 ) )   n = 22   d_n = 1+1i 
assign Y[4'b0101] [23] = 144'h 000000000000000001000000000008000000;  // 000000000FFFFFE000 +0.0000001192092753 =  1 * atan( 1 / (  1 + 2^23 ) )   n = 23   d_n = 1+1i 
assign Y[4'b0101] [24] = 144'h 000000000000000000400000000000800000;  // 0000000007FFFFF800 +0.0000000596046412 =  1 * atan( 1 / (  1 + 2^24 ) )   n = 24   d_n = 1+1i 
assign Y[4'b0101] [25] = 144'h 000000000000000000100000000000080000;  // 0000000003FFFFFE00 +0.0000000298023215 =  1 * atan( 1 / (  1 + 2^25 ) )   n = 25   d_n = 1+1i 
assign Y[4'b0101] [26] = 144'h 000000000000000000040000000000008000;  // 0000000001FFFFFF80 +0.0000000149011610 =  1 * atan( 1 / (  1 + 2^26 ) )   n = 26   d_n = 1+1i 
assign Y[4'b0101] [27] = 144'h 000000000000000000010000000000000800;  // 0000000000FFFFFFE0 +0.0000000074505805 =  1 * atan( 1 / (  1 + 2^27 ) )   n = 27   d_n = 1+1i 
assign Y[4'b0101] [28] = 144'h 000000000000000000004000000000000080;  // 00000000007FFFFFF8 +0.0000000037252903 =  1 * atan( 1 / (  1 + 2^28 ) )   n = 28   d_n = 1+1i 
assign Y[4'b0101] [29] = 144'h 000000000000000000001000000000000008;  // 00000000003FFFFFFE +0.0000000018626451 =  1 * atan( 1 / (  1 + 2^29 ) )   n = 29   d_n = 1+1i 
assign Y[4'b0101] [30] = 144'h 000000000000000000000400000000000000;  // 00000000001FFFFFFF +0.0000000009313226 =  1 * atan( 1 / (  1 + 2^30 ) )   n = 30   d_n = 1+1i 
assign Y[4'b0101] [31] = 144'h 000000000000000000000100000000000000;  // 00000000000FFFFFFF +0.0000000004656613 =  1 * atan( 1 / (  1 + 2^31 ) )   n = 31   d_n = 1+1i 
assign Y[4'b0101] [32] = 144'h 000000000000000000000040000000000000;  // 000000000007FFFFFF +0.0000000002328306 =  1 * atan( 1 / (  1 + 2^32 ) )   n = 32   d_n = 1+1i 
assign Y[4'b0101] [33] = 144'h 000000000000000000000010000000000000;  // 000000000003FFFFFF +0.0000000001164153 =  1 * atan( 1 / (  1 + 2^33 ) )   n = 33   d_n = 1+1i 
assign Y[4'b0101] [34] = 144'h 000000000000000000000004000000000000;  // 000000000001FFFFFF +0.0000000000582077 =  1 * atan( 1 / (  1 + 2^34 ) )   n = 34   d_n = 1+1i 
assign Y[4'b0101] [35] = 144'h 000000000000000000000001000000000000;  // 000000000000FFFFFF +0.0000000000291038 =  1 * atan( 1 / (  1 + 2^35 ) )   n = 35   d_n = 1+1i 
assign Y[4'b0101] [36] = 144'h 000000000000000000000000400000000000;  // 0000000000007FFFFF +0.0000000000145519 =  1 * atan( 1 / (  1 + 2^36 ) )   n = 36   d_n = 1+1i 
assign Y[4'b0101] [37] = 144'h 000000000000000000000000100000000000;  // 0000000000003FFFFF +0.0000000000072760 =  1 * atan( 1 / (  1 + 2^37 ) )   n = 37   d_n = 1+1i 
assign Y[4'b0101] [38] = 144'h 000000000000000000000000040000000000;  // 0000000000001FFFFF +0.0000000000036380 =  1 * atan( 1 / (  1 + 2^38 ) )   n = 38   d_n = 1+1i 
assign Y[4'b0101] [39] = 144'h 000000000000000000000000010000000000;  // 0000000000000FFFFF +0.0000000000018190 =  1 * atan( 1 / (  1 + 2^39 ) )   n = 39   d_n = 1+1i 
assign Y[4'b0101] [40] = 144'h 000000000000000000000000004000000000;  // 00000000000007FFFF +0.0000000000009095 =  1 * atan( 1 / (  1 + 2^40 ) )   n = 40   d_n = 1+1i 
assign Y[4'b0101] [41] = 144'h 000000000000000000000000001000000000;  // 00000000000003FFFF +0.0000000000004547 =  1 * atan( 1 / (  1 + 2^41 ) )   n = 41   d_n = 1+1i 
assign Y[4'b0101] [42] = 144'h 000000000000000000000000000400000000;  // 00000000000001FFFF +0.0000000000002274 =  1 * atan( 1 / (  1 + 2^42 ) )   n = 42   d_n = 1+1i 
assign Y[4'b0101] [43] = 144'h 000000000000000000000000000100000000;  // 00000000000000FFFF +0.0000000000001137 =  1 * atan( 1 / (  1 + 2^43 ) )   n = 43   d_n = 1+1i 
assign Y[4'b0101] [44] = 144'h 000000000000000000000000000040000000;  // 000000000000007FFF +0.0000000000000568 =  1 * atan( 1 / (  1 + 2^44 ) )   n = 44   d_n = 1+1i 
assign Y[4'b0101] [45] = 144'h 000000000000000000000000000010000000;  // 000000000000003FFF +0.0000000000000284 =  1 * atan( 1 / (  1 + 2^45 ) )   n = 45   d_n = 1+1i 
assign Y[4'b0101] [46] = 144'h 000000000000000000000000000004000000;  // 000000000000001FFF +0.0000000000000142 =  1 * atan( 1 / (  1 + 2^46 ) )   n = 46   d_n = 1+1i 
assign Y[4'b0101] [47] = 144'h 000000000000000000000000000001000000;  // 000000000000000FFF +0.0000000000000071 =  1 * atan( 1 / (  1 + 2^47 ) )   n = 47   d_n = 1+1i 
assign Y[4'b0101] [48] = 144'h 000000000000000000000000000000400000;  // 0000000000000007FF +0.0000000000000036 =  1 * atan( 1 / (  1 + 2^48 ) )   n = 48   d_n = 1+1i 
assign Y[4'b0101] [49] = 144'h 000000000000000000000000000000100000;  // 0000000000000003FF +0.0000000000000018 =  1 * atan( 1 / (  1 + 2^49 ) )   n = 49   d_n = 1+1i 
assign Y[4'b0101] [50] = 144'h 000000000000000000000000000000040000;  // 0000000000000001FF +0.0000000000000009 =  1 * atan( 1 / (  1 + 2^50 ) )   n = 50   d_n = 1+1i 
assign Y[4'b0101] [51] = 144'h 000000000000000000000000000000010000;  // 0000000000000000FF +0.0000000000000004 =  1 * atan( 1 / (  1 + 2^51 ) )   n = 51   d_n = 1+1i 
assign Y[4'b0101] [52] = 144'h 000000000000000000000000000000004000;  // 00000000000000007F +0.0000000000000002 =  1 * atan( 1 / (  1 + 2^52 ) )   n = 52   d_n = 1+1i 
assign Y[4'b0101] [53] = 144'h 000000000000000000000000000000001000;  // 000000000000000040 +0.0000000000000001 =  1 * atan( 1 / (  1 + 2^53 ) )   n = 53   d_n = 1+1i 
assign Y[4'b0101] [54] = 144'h 000000000000000000000000000000000400;  // 000000000000000020 +0.0000000000000001 =  1 * atan( 1 / (  1 + 2^54 ) )   n = 54   d_n = 1+1i 
assign Y[4'b0101] [55] = 144'h 000000000000000000000000000000000100;  // 000000000000000010 +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^55 ) )   n = 55   d_n = 1+1i 
assign Y[4'b0101] [56] = 144'h 000000000000000000000000000000000040;  // 000000000000000008 +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^56 ) )   n = 56   d_n = 1+1i 
assign Y[4'b0101] [57] = 144'h 000000000000000000000000000000000010;  // 000000000000000004 +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^57 ) )   n = 57   d_n = 1+1i 
assign Y[4'b0101] [58] = 144'h 000000000000000000000000000000000004;  // 000000000000000002 +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^58 ) )   n = 58   d_n = 1+1i 
assign Y[4'b0101] [59] = 144'h 000000000000000000000000000000000001;  // 000000000000000001 +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^59 ) )   n = 59   d_n = 1+1i 
assign Y[4'b0101] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^60 ) )   n = 60   d_n = 1+1i 
assign Y[4'b0101] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^61 ) )   n = 61   d_n = 1+1i 
assign Y[4'b0101] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^62 ) )   n = 62   d_n = 1+1i 
assign Y[4'b0101] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^63 ) )   n = 63   d_n = 1+1i 
assign Y[4'b0101] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / (  1 + 2^64 ) )   n = 64   d_n = 1+1i 
assign Y[4'b0110] [01] = 144'h 000000102088812108012220108088440800;  // 0003B58CE0AC3769E0 +0.4636476090008061 =  1 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = 0+1i 
assign Y[4'b0110] [02] = 144'h 000000040088208088008112204001082000;  // 0001F5B75F92C80DD0 +0.2449786631268641 =  1 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = 0+1i 
assign Y[4'b0110] [03] = 144'h 000000010002220821110888880480208200;  // 0000FEADD4D5617B70 +0.1243549945467614 =  1 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = 0+1i 
assign Y[4'b0110] [04] = 144'h 000000004000088882020821221000808440;  // 00007FD56EDCB3F7A8 +0.0624188099959574 =  1 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = 0+1i 
assign Y[4'b0110] [05] = 144'h 000000001000002222208082111202201040;  // 00003FFAAB7752EC4A +0.0312398334302683 =  1 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = 0+1i 
assign Y[4'b0110] [06] = 144'h 000000000400000088888820202082044422;  // 00001FFF555BBB729B +0.0156237286204768 =  1 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = 0+1i 
assign Y[4'b0110] [07] = 144'h 000000000100000002222222080808211120;  // 00000FFFEAAADDDD4B +0.0078123410601011 =  1 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = 0+1i 
assign Y[4'b0110] [08] = 144'h 000000000040000000088888888202020208;  // 000007FFFD5556EEED +0.0039062301319670 =  1 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = 0+1i 
assign Y[4'b0110] [09] = 144'h 000000000010000000002222222220808080;  // 000003FFFFAAAAB777 +0.0019531225164788 =  1 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = 0+1i 
assign Y[4'b0110] [10] = 144'h 000000000004000000000088888888882020;  // 000001FFFFF55555BB +0.0009765621895593 =  1 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = 0+1i 
assign Y[4'b0110] [11] = 144'h 000000000001000000000002222222222208;  // 000000FFFFFEAAAAAD +0.0004882812111949 =  1 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = 0+1i 
assign Y[4'b0110] [12] = 144'h 000000000000400000000000088888888888;  // 0000007FFFFFD55555 +0.0002441406201494 =  1 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = 0+1i 
assign Y[4'b0110] [13] = 144'h 000000000000100000000000008444444444;  // 0000003FFFFFFAAAAA +0.0001220703118937 =  1 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = 0+1i 
assign Y[4'b0110] [14] = 144'h 000000000000040000000000000211111111;  // 0000001FFFFFFF5555 +0.0000610351561742 =  1 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = 0+1i 
assign Y[4'b0110] [15] = 144'h 000000000000010000000000000008444444;  // 0000000FFFFFFFEAAA +0.0000305175781155 =  1 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = 0+1i 
assign Y[4'b0110] [16] = 144'h 000000000000004000000000000000211111;  // 00000007FFFFFFFD55 +0.0000152587890613 =  1 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = 0+1i 
assign Y[4'b0110] [17] = 144'h 000000000000001000000000000000008444;  // 00000003FFFFFFFFAA +0.0000076293945311 =  1 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = 0+1i 
assign Y[4'b0110] [18] = 144'h 000000000000000400000000000000000211;  // 00000001FFFFFFFFF5 +0.0000038146972656 =  1 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = 0+1i 
assign Y[4'b0110] [19] = 144'h 000000000000000100000000000000000008;  // 00000000FFFFFFFFFE +0.0000019073486328 =  1 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = 0+1i 
assign Y[4'b0110] [20] = 144'h 000000000000000040000000000000000000;  // 000000007FFFFFFFFF +0.0000009536743164 =  1 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = 0+1i 
assign Y[4'b0110] [21] = 144'h 000000000000000010000000000000000000;  // 000000003FFFFFFFFF +0.0000004768371582 =  1 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = 0+1i 
assign Y[4'b0110] [22] = 144'h 000000000000000004000000000000000000;  // 000000001FFFFFFFFF +0.0000002384185791 =  1 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = 0+1i 
assign Y[4'b0110] [23] = 144'h 000000000000000001000000000000000000;  // 000000000FFFFFFFFF +0.0000001192092896 =  1 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = 0+1i 
assign Y[4'b0110] [24] = 144'h 000000000000000000400000000000000000;  // 0000000007FFFFFFFF +0.0000000596046448 =  1 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = 0+1i 
assign Y[4'b0110] [25] = 144'h 000000000000000000100000000000000000;  // 0000000003FFFFFFFF +0.0000000298023224 =  1 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = 0+1i 
assign Y[4'b0110] [26] = 144'h 000000000000000000040000000000000000;  // 0000000001FFFFFFFF +0.0000000149011612 =  1 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = 0+1i 
assign Y[4'b0110] [27] = 144'h 000000000000000000010000000000000000;  // 000000000100000000 +0.0000000074505806 =  1 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = 0+1i 
assign Y[4'b0110] [28] = 144'h 000000000000000000004000000000000000;  // 000000000080000000 +0.0000000037252903 =  1 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = 0+1i 
assign Y[4'b0110] [29] = 144'h 000000000000000000001000000000000000;  // 000000000040000000 +0.0000000018626451 =  1 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = 0+1i 
assign Y[4'b0110] [30] = 144'h 000000000000000000000400000000000000;  // 000000000020000000 +0.0000000009313226 =  1 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = 0+1i 
assign Y[4'b0110] [31] = 144'h 000000000000000000000100000000000000;  // 000000000010000000 +0.0000000004656613 =  1 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = 0+1i 
assign Y[4'b0110] [32] = 144'h 000000000000000000000040000000000000;  // 000000000008000000 +0.0000000002328306 =  1 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = 0+1i 
assign Y[4'b0110] [33] = 144'h 000000000000000000000010000000000000;  // 000000000004000000 +0.0000000001164153 =  1 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = 0+1i 
assign Y[4'b0110] [34] = 144'h 000000000000000000000004000000000000;  // 000000000002000000 +0.0000000000582077 =  1 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = 0+1i 
assign Y[4'b0110] [35] = 144'h 000000000000000000000001000000000000;  // 000000000001000000 +0.0000000000291038 =  1 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = 0+1i 
assign Y[4'b0110] [36] = 144'h 000000000000000000000000400000000000;  // 000000000000800000 +0.0000000000145519 =  1 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = 0+1i 
assign Y[4'b0110] [37] = 144'h 000000000000000000000000100000000000;  // 000000000000400000 +0.0000000000072760 =  1 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = 0+1i 
assign Y[4'b0110] [38] = 144'h 000000000000000000000000040000000000;  // 000000000000200000 +0.0000000000036380 =  1 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = 0+1i 
assign Y[4'b0110] [39] = 144'h 000000000000000000000000010000000000;  // 000000000000100000 +0.0000000000018190 =  1 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = 0+1i 
assign Y[4'b0110] [40] = 144'h 000000000000000000000000004000000000;  // 000000000000080000 +0.0000000000009095 =  1 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = 0+1i 
assign Y[4'b0110] [41] = 144'h 000000000000000000000000001000000000;  // 000000000000040000 +0.0000000000004547 =  1 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = 0+1i 
assign Y[4'b0110] [42] = 144'h 000000000000000000000000000400000000;  // 000000000000020000 +0.0000000000002274 =  1 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = 0+1i 
assign Y[4'b0110] [43] = 144'h 000000000000000000000000000100000000;  // 000000000000010000 +0.0000000000001137 =  1 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = 0+1i 
assign Y[4'b0110] [44] = 144'h 000000000000000000000000000040000000;  // 000000000000008000 +0.0000000000000568 =  1 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = 0+1i 
assign Y[4'b0110] [45] = 144'h 000000000000000000000000000010000000;  // 000000000000004000 +0.0000000000000284 =  1 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = 0+1i 
assign Y[4'b0110] [46] = 144'h 000000000000000000000000000004000000;  // 000000000000002000 +0.0000000000000142 =  1 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = 0+1i 
assign Y[4'b0110] [47] = 144'h 000000000000000000000000000001000000;  // 000000000000001000 +0.0000000000000071 =  1 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = 0+1i 
assign Y[4'b0110] [48] = 144'h 000000000000000000000000000000400000;  // 000000000000000800 +0.0000000000000036 =  1 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = 0+1i 
assign Y[4'b0110] [49] = 144'h 000000000000000000000000000000100000;  // 000000000000000400 +0.0000000000000018 =  1 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = 0+1i 
assign Y[4'b0110] [50] = 144'h 000000000000000000000000000000040000;  // 000000000000000200 +0.0000000000000009 =  1 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = 0+1i 
assign Y[4'b0110] [51] = 144'h 000000000000000000000000000000010000;  // 000000000000000100 +0.0000000000000004 =  1 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = 0+1i 
assign Y[4'b0110] [52] = 144'h 000000000000000000000000000000004000;  // 000000000000000080 +0.0000000000000002 =  1 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = 0+1i 
assign Y[4'b0110] [53] = 144'h 000000000000000000000000000000001000;  // 000000000000000040 +0.0000000000000001 =  1 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = 0+1i 
assign Y[4'b0110] [54] = 144'h 000000000000000000000000000000000400;  // 000000000000000020 +0.0000000000000001 =  1 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = 0+1i 
assign Y[4'b0110] [55] = 144'h 000000000000000000000000000000000100;  // 000000000000000010 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = 0+1i 
assign Y[4'b0110] [56] = 144'h 000000000000000000000000000000000040;  // 000000000000000008 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = 0+1i 
assign Y[4'b0110] [57] = 144'h 000000000000000000000000000000000010;  // 000000000000000004 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = 0+1i 
assign Y[4'b0110] [58] = 144'h 000000000000000000000000000000000004;  // 000000000000000002 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = 0+1i 
assign Y[4'b0110] [59] = 144'h 000000000000000000000000000000000001;  // 000000000000000001 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = 0+1i 
assign Y[4'b0110] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = 0+1i 
assign Y[4'b0110] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = 0+1i 
assign Y[4'b0110] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = 0+1i 
assign Y[4'b0110] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = 0+1i 
assign Y[4'b0110] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = 0+1i 
assign Y[4'b0111] [01] = 144'h 000000481040400221110101012210480000;  // 0006487ED5110B4600 +0.7853981633974483 =  1 * atan( 1 / ( -1 + 2^1 ) )   n =  1   d_n = -1+1i 
assign Y[4'b0111] [02] = 144'h 000000044112020402104811211008200400;  // 000292F1F464D3DC20 +0.3217505543966422 =  1 * atan( 1 / ( -1 + 2^2 ) )   n =  2   d_n = -1+1i 
assign Y[4'b0111] [03] = 144'h 000000010404442202201040881081082100;  // 0001229AEC47638DD0 +0.1418970546041639 =  1 * atan( 1 / ( -1 + 2^3 ) )   n =  3   d_n = -1+1i 
assign Y[4'b0111] [04] = 144'h 000000004040111108102212008420810400;  // 00008854E3B2F9B920 +0.0665681637758238 =  1 * atan( 1 / ( -1 + 2^4 ) )   n =  4   d_n = -1+1i 
assign Y[4'b0111] [05] = 144'h 000000001004004444421120844122120800;  // 0000420AA74BA8B2E0 +0.0322468824352539 =  1 * atan( 1 / ( -1 + 2^5 ) )   n =  5   d_n = -1+1i 
assign Y[4'b0111] [06] = 144'h 000000000400400111111022010220400440;  // 00002081553B0EC828 +0.0158716829917901 =  1 * atan( 1 / ( -1 + 2^6 ) )   n =  6   d_n = -1+1i 
assign Y[4'b0111] [07] = 144'h 000000000100040004444444082212084401;  // 000010202AA9DB2EA1 +0.0078738530241005 =  1 * atan( 1 / ( -1 + 2^7 ) )   n =  7   d_n = -1+1i 
assign Y[4'b0111] [08] = 144'h 000000000040004000111111110208101022;  // 0000080805554EE43B +0.0039215485247600 =  1 * atan( 1 / ( -1 + 2^8 ) )   n =  8   d_n = -1+1i 
assign Y[4'b0111] [09] = 144'h 000000000010000400004444444440821121;  // 0000040200AAAA774C +0.0019569446642965 =  1 * atan( 1 / ( -1 + 2^9 ) )   n =  9   d_n = -1+1i 
assign Y[4'b0111] [10] = 144'h 000000000004000040000111111111102022;  // 0000020080155553BB +0.0009775167951974 =  1 * atan( 1 / ( -1 + 2^10 ) )   n = 10   d_n = -1+1i 
assign Y[4'b0111] [11] = 144'h 000000000001000004000004444444444408;  // 000001002002AAAA9D +0.0004885197461893 =  1 * atan( 1 / ( -1 + 2^11 ) )   n = 11   d_n = -1+1i 
assign Y[4'b0111] [12] = 144'h 000000000000400000400000111111111111;  // 000000800800555554 +0.0002442002393461 =  1 * atan( 1 / ( -1 + 2^12 ) )   n = 12   d_n = -1+1i 
assign Y[4'b0111] [13] = 144'h 000000000000100000040000004444444444;  // 0000004002000AAAAA +0.0001220852148739 =  1 * atan( 1 / ( -1 + 2^13 ) )   n = 13   d_n = -1+1i 
assign Y[4'b0111] [14] = 144'h 000000000000040000004000000111111111;  // 000000200080015555 +0.0000610388816919 =  1 * atan( 1 / ( -1 + 2^14 ) )   n = 14   d_n = -1+1i 
assign Y[4'b0111] [15] = 144'h 000000000000010000000400000004444444;  // 000000100020002AAA +0.0000305185094665 =  1 * atan( 1 / ( -1 + 2^15 ) )   n = 15   d_n = -1+1i 
assign Y[4'b0111] [16] = 144'h 000000000000004000000040000000111111;  // 000000080008000555 +0.0000152590218955 =  1 * atan( 1 / ( -1 + 2^16 ) )   n = 16   d_n = -1+1i 
assign Y[4'b0111] [17] = 144'h 000000000000001000000004000000004444;  // 0000000400020000AA +0.0000076294527392 =  1 * atan( 1 / ( -1 + 2^17 ) )   n = 17   d_n = -1+1i 
assign Y[4'b0111] [18] = 144'h 000000000000000400000000400000000111;  // 000000020000800015 +0.0000038147118176 =  1 * atan( 1 / ( -1 + 2^18 ) )   n = 18   d_n = -1+1i 
assign Y[4'b0111] [19] = 144'h 000000000000000100000000040000000004;  // 000000010000200002 +0.0000019073522708 =  1 * atan( 1 / ( -1 + 2^19 ) )   n = 19   d_n = -1+1i 
assign Y[4'b0111] [20] = 144'h 000000000000000040000000004000000000;  // 000000008000080000 +0.0000009536752259 =  1 * atan( 1 / ( -1 + 2^20 ) )   n = 20   d_n = -1+1i 
assign Y[4'b0111] [21] = 144'h 000000000000000010000000000400000000;  // 000000004000020000 +0.0000004768373856 =  1 * atan( 1 / ( -1 + 2^21 ) )   n = 21   d_n = -1+1i 
assign Y[4'b0111] [22] = 144'h 000000000000000004000000000040000000;  // 000000002000008000 +0.0000002384186359 =  1 * atan( 1 / ( -1 + 2^22 ) )   n = 22   d_n = -1+1i 
assign Y[4'b0111] [23] = 144'h 000000000000000001000000000004000000;  // 000000001000002000 +0.0000001192093038 =  1 * atan( 1 / ( -1 + 2^23 ) )   n = 23   d_n = -1+1i 
assign Y[4'b0111] [24] = 144'h 000000000000000000400000000000400000;  // 000000000800000800 +0.0000000596046483 =  1 * atan( 1 / ( -1 + 2^24 ) )   n = 24   d_n = -1+1i 
assign Y[4'b0111] [25] = 144'h 000000000000000000100000000000040000;  // 000000000400000200 +0.0000000298023233 =  1 * atan( 1 / ( -1 + 2^25 ) )   n = 25   d_n = -1+1i 
assign Y[4'b0111] [26] = 144'h 000000000000000000040000000000004000;  // 000000000200000080 +0.0000000149011614 =  1 * atan( 1 / ( -1 + 2^26 ) )   n = 26   d_n = -1+1i 
assign Y[4'b0111] [27] = 144'h 000000000000000000010000000000000400;  // 000000000100000020 +0.0000000074505807 =  1 * atan( 1 / ( -1 + 2^27 ) )   n = 27   d_n = -1+1i 
assign Y[4'b0111] [28] = 144'h 000000000000000000004000000000000040;  // 000000000080000008 +0.0000000037252903 =  1 * atan( 1 / ( -1 + 2^28 ) )   n = 28   d_n = -1+1i 
assign Y[4'b0111] [29] = 144'h 000000000000000000001000000000000004;  // 000000000040000002 +0.0000000018626452 =  1 * atan( 1 / ( -1 + 2^29 ) )   n = 29   d_n = -1+1i 
assign Y[4'b0111] [30] = 144'h 000000000000000000000400000000000000;  // 000000000020000000 +0.0000000009313226 =  1 * atan( 1 / ( -1 + 2^30 ) )   n = 30   d_n = -1+1i 
assign Y[4'b0111] [31] = 144'h 000000000000000000000100000000000000;  // 000000000010000000 +0.0000000004656613 =  1 * atan( 1 / ( -1 + 2^31 ) )   n = 31   d_n = -1+1i 
assign Y[4'b0111] [32] = 144'h 000000000000000000000040000000000000;  // 000000000008000000 +0.0000000002328306 =  1 * atan( 1 / ( -1 + 2^32 ) )   n = 32   d_n = -1+1i 
assign Y[4'b0111] [33] = 144'h 000000000000000000000010000000000000;  // 000000000004000000 +0.0000000001164153 =  1 * atan( 1 / ( -1 + 2^33 ) )   n = 33   d_n = -1+1i 
assign Y[4'b0111] [34] = 144'h 000000000000000000000004000000000000;  // 000000000002000000 +0.0000000000582077 =  1 * atan( 1 / ( -1 + 2^34 ) )   n = 34   d_n = -1+1i 
assign Y[4'b0111] [35] = 144'h 000000000000000000000001000000000000;  // 000000000001000000 +0.0000000000291038 =  1 * atan( 1 / ( -1 + 2^35 ) )   n = 35   d_n = -1+1i 
assign Y[4'b0111] [36] = 144'h 000000000000000000000000400000000000;  // 000000000000800000 +0.0000000000145519 =  1 * atan( 1 / ( -1 + 2^36 ) )   n = 36   d_n = -1+1i 
assign Y[4'b0111] [37] = 144'h 000000000000000000000000100000000000;  // 000000000000400000 +0.0000000000072760 =  1 * atan( 1 / ( -1 + 2^37 ) )   n = 37   d_n = -1+1i 
assign Y[4'b0111] [38] = 144'h 000000000000000000000000040000000000;  // 000000000000200000 +0.0000000000036380 =  1 * atan( 1 / ( -1 + 2^38 ) )   n = 38   d_n = -1+1i 
assign Y[4'b0111] [39] = 144'h 000000000000000000000000010000000000;  // 000000000000100000 +0.0000000000018190 =  1 * atan( 1 / ( -1 + 2^39 ) )   n = 39   d_n = -1+1i 
assign Y[4'b0111] [40] = 144'h 000000000000000000000000004000000000;  // 000000000000080000 +0.0000000000009095 =  1 * atan( 1 / ( -1 + 2^40 ) )   n = 40   d_n = -1+1i 
assign Y[4'b0111] [41] = 144'h 000000000000000000000000001000000000;  // 000000000000040000 +0.0000000000004547 =  1 * atan( 1 / ( -1 + 2^41 ) )   n = 41   d_n = -1+1i 
assign Y[4'b0111] [42] = 144'h 000000000000000000000000000400000000;  // 000000000000020000 +0.0000000000002274 =  1 * atan( 1 / ( -1 + 2^42 ) )   n = 42   d_n = -1+1i 
assign Y[4'b0111] [43] = 144'h 000000000000000000000000000100000000;  // 000000000000010000 +0.0000000000001137 =  1 * atan( 1 / ( -1 + 2^43 ) )   n = 43   d_n = -1+1i 
assign Y[4'b0111] [44] = 144'h 000000000000000000000000000040000000;  // 000000000000008000 +0.0000000000000568 =  1 * atan( 1 / ( -1 + 2^44 ) )   n = 44   d_n = -1+1i 
assign Y[4'b0111] [45] = 144'h 000000000000000000000000000010000000;  // 000000000000004000 +0.0000000000000284 =  1 * atan( 1 / ( -1 + 2^45 ) )   n = 45   d_n = -1+1i 
assign Y[4'b0111] [46] = 144'h 000000000000000000000000000004000000;  // 000000000000002000 +0.0000000000000142 =  1 * atan( 1 / ( -1 + 2^46 ) )   n = 46   d_n = -1+1i 
assign Y[4'b0111] [47] = 144'h 000000000000000000000000000001000000;  // 000000000000001000 +0.0000000000000071 =  1 * atan( 1 / ( -1 + 2^47 ) )   n = 47   d_n = -1+1i 
assign Y[4'b0111] [48] = 144'h 000000000000000000000000000000400000;  // 000000000000000800 +0.0000000000000036 =  1 * atan( 1 / ( -1 + 2^48 ) )   n = 48   d_n = -1+1i 
assign Y[4'b0111] [49] = 144'h 000000000000000000000000000000100000;  // 000000000000000400 +0.0000000000000018 =  1 * atan( 1 / ( -1 + 2^49 ) )   n = 49   d_n = -1+1i 
assign Y[4'b0111] [50] = 144'h 000000000000000000000000000000040000;  // 000000000000000200 +0.0000000000000009 =  1 * atan( 1 / ( -1 + 2^50 ) )   n = 50   d_n = -1+1i 
assign Y[4'b0111] [51] = 144'h 000000000000000000000000000000010000;  // 000000000000000100 +0.0000000000000004 =  1 * atan( 1 / ( -1 + 2^51 ) )   n = 51   d_n = -1+1i 
assign Y[4'b0111] [52] = 144'h 000000000000000000000000000000004000;  // 000000000000000080 +0.0000000000000002 =  1 * atan( 1 / ( -1 + 2^52 ) )   n = 52   d_n = -1+1i 
assign Y[4'b0111] [53] = 144'h 000000000000000000000000000000001000;  // 000000000000000040 +0.0000000000000001 =  1 * atan( 1 / ( -1 + 2^53 ) )   n = 53   d_n = -1+1i 
assign Y[4'b0111] [54] = 144'h 000000000000000000000000000000000400;  // 000000000000000020 +0.0000000000000001 =  1 * atan( 1 / ( -1 + 2^54 ) )   n = 54   d_n = -1+1i 
assign Y[4'b0111] [55] = 144'h 000000000000000000000000000000000100;  // 000000000000000010 +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^55 ) )   n = 55   d_n = -1+1i 
assign Y[4'b0111] [56] = 144'h 000000000000000000000000000000000040;  // 000000000000000008 +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^56 ) )   n = 56   d_n = -1+1i 
assign Y[4'b0111] [57] = 144'h 000000000000000000000000000000000010;  // 000000000000000004 +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^57 ) )   n = 57   d_n = -1+1i 
assign Y[4'b0111] [58] = 144'h 000000000000000000000000000000000004;  // 000000000000000002 +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^58 ) )   n = 58   d_n = -1+1i 
assign Y[4'b0111] [59] = 144'h 000000000000000000000000000000000001;  // 000000000000000001 +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^59 ) )   n = 59   d_n = -1+1i 
assign Y[4'b0111] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^60 ) )   n = 60   d_n = -1+1i 
assign Y[4'b0111] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^61 ) )   n = 61   d_n = -1+1i 
assign Y[4'b0111] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^62 ) )   n = 62   d_n = -1+1i 
assign Y[4'b0111] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^63 ) )   n = 63   d_n = -1+1i 
assign Y[4'b0111] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  1 * atan( 1 / ( -1 + 2^64 ) )   n = 64   d_n = -1+1i 
assign Y[4'b1000] [01] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = 0 
assign Y[4'b1000] [02] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = 0 
assign Y[4'b1000] [03] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = 0 
assign Y[4'b1000] [04] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = 0 
assign Y[4'b1000] [05] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = 0 
assign Y[4'b1000] [06] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = 0 
assign Y[4'b1000] [07] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = 0 
assign Y[4'b1000] [08] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = 0 
assign Y[4'b1000] [09] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = 0 
assign Y[4'b1000] [10] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = 0 
assign Y[4'b1000] [11] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = 0 
assign Y[4'b1000] [12] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = 0 
assign Y[4'b1000] [13] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = 0 
assign Y[4'b1000] [14] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = 0 
assign Y[4'b1000] [15] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = 0 
assign Y[4'b1000] [16] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = 0 
assign Y[4'b1000] [17] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = 0 
assign Y[4'b1000] [18] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = 0 
assign Y[4'b1000] [19] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = 0 
assign Y[4'b1000] [20] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = 0 
assign Y[4'b1000] [21] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = 0 
assign Y[4'b1000] [22] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = 0 
assign Y[4'b1000] [23] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = 0 
assign Y[4'b1000] [24] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = 0 
assign Y[4'b1000] [25] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = 0 
assign Y[4'b1000] [26] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = 0 
assign Y[4'b1000] [27] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = 0 
assign Y[4'b1000] [28] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = 0 
assign Y[4'b1000] [29] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = 0 
assign Y[4'b1000] [30] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = 0 
assign Y[4'b1000] [31] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = 0 
assign Y[4'b1000] [32] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = 0 
assign Y[4'b1000] [33] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = 0 
assign Y[4'b1000] [34] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = 0 
assign Y[4'b1000] [35] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = 0 
assign Y[4'b1000] [36] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = 0 
assign Y[4'b1000] [37] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = 0 
assign Y[4'b1000] [38] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = 0 
assign Y[4'b1000] [39] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = 0 
assign Y[4'b1000] [40] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = 0 
assign Y[4'b1000] [41] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = 0 
assign Y[4'b1000] [42] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = 0 
assign Y[4'b1000] [43] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = 0 
assign Y[4'b1000] [44] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = 0 
assign Y[4'b1000] [45] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = 0 
assign Y[4'b1000] [46] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = 0 
assign Y[4'b1000] [47] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = 0 
assign Y[4'b1000] [48] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = 0 
assign Y[4'b1000] [49] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = 0 
assign Y[4'b1000] [50] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = 0 
assign Y[4'b1000] [51] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = 0 
assign Y[4'b1000] [52] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = 0 
assign Y[4'b1000] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = 0 
assign Y[4'b1000] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = 0 
assign Y[4'b1000] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = 0 
assign Y[4'b1000] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = 0 
assign Y[4'b1000] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = 0 
assign Y[4'b1000] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = 0 
assign Y[4'b1000] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = 0 
assign Y[4'b1000] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = 0 
assign Y[4'b1000] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = 0 
assign Y[4'b1000] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = 0 
assign Y[4'b1000] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = 0 
assign Y[4'b1000] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = 0 
assign Y[4'b1001] [01] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^1 ) )   n =  1   d_n = 1 
assign Y[4'b1001] [02] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^2 ) )   n =  2   d_n = 1 
assign Y[4'b1001] [03] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^3 ) )   n =  3   d_n = 1 
assign Y[4'b1001] [04] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^4 ) )   n =  4   d_n = 1 
assign Y[4'b1001] [05] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^5 ) )   n =  5   d_n = 1 
assign Y[4'b1001] [06] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^6 ) )   n =  6   d_n = 1 
assign Y[4'b1001] [07] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^7 ) )   n =  7   d_n = 1 
assign Y[4'b1001] [08] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^8 ) )   n =  8   d_n = 1 
assign Y[4'b1001] [09] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^9 ) )   n =  9   d_n = 1 
assign Y[4'b1001] [10] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^10 ) )   n = 10   d_n = 1 
assign Y[4'b1001] [11] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^11 ) )   n = 11   d_n = 1 
assign Y[4'b1001] [12] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^12 ) )   n = 12   d_n = 1 
assign Y[4'b1001] [13] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^13 ) )   n = 13   d_n = 1 
assign Y[4'b1001] [14] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^14 ) )   n = 14   d_n = 1 
assign Y[4'b1001] [15] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^15 ) )   n = 15   d_n = 1 
assign Y[4'b1001] [16] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^16 ) )   n = 16   d_n = 1 
assign Y[4'b1001] [17] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^17 ) )   n = 17   d_n = 1 
assign Y[4'b1001] [18] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^18 ) )   n = 18   d_n = 1 
assign Y[4'b1001] [19] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^19 ) )   n = 19   d_n = 1 
assign Y[4'b1001] [20] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^20 ) )   n = 20   d_n = 1 
assign Y[4'b1001] [21] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^21 ) )   n = 21   d_n = 1 
assign Y[4'b1001] [22] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^22 ) )   n = 22   d_n = 1 
assign Y[4'b1001] [23] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^23 ) )   n = 23   d_n = 1 
assign Y[4'b1001] [24] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^24 ) )   n = 24   d_n = 1 
assign Y[4'b1001] [25] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^25 ) )   n = 25   d_n = 1 
assign Y[4'b1001] [26] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^26 ) )   n = 26   d_n = 1 
assign Y[4'b1001] [27] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^27 ) )   n = 27   d_n = 1 
assign Y[4'b1001] [28] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^28 ) )   n = 28   d_n = 1 
assign Y[4'b1001] [29] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^29 ) )   n = 29   d_n = 1 
assign Y[4'b1001] [30] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^30 ) )   n = 30   d_n = 1 
assign Y[4'b1001] [31] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^31 ) )   n = 31   d_n = 1 
assign Y[4'b1001] [32] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^32 ) )   n = 32   d_n = 1 
assign Y[4'b1001] [33] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^33 ) )   n = 33   d_n = 1 
assign Y[4'b1001] [34] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^34 ) )   n = 34   d_n = 1 
assign Y[4'b1001] [35] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^35 ) )   n = 35   d_n = 1 
assign Y[4'b1001] [36] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^36 ) )   n = 36   d_n = 1 
assign Y[4'b1001] [37] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^37 ) )   n = 37   d_n = 1 
assign Y[4'b1001] [38] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^38 ) )   n = 38   d_n = 1 
assign Y[4'b1001] [39] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^39 ) )   n = 39   d_n = 1 
assign Y[4'b1001] [40] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^40 ) )   n = 40   d_n = 1 
assign Y[4'b1001] [41] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^41 ) )   n = 41   d_n = 1 
assign Y[4'b1001] [42] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^42 ) )   n = 42   d_n = 1 
assign Y[4'b1001] [43] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^43 ) )   n = 43   d_n = 1 
assign Y[4'b1001] [44] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^44 ) )   n = 44   d_n = 1 
assign Y[4'b1001] [45] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^45 ) )   n = 45   d_n = 1 
assign Y[4'b1001] [46] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^46 ) )   n = 46   d_n = 1 
assign Y[4'b1001] [47] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^47 ) )   n = 47   d_n = 1 
assign Y[4'b1001] [48] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^48 ) )   n = 48   d_n = 1 
assign Y[4'b1001] [49] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^49 ) )   n = 49   d_n = 1 
assign Y[4'b1001] [50] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^50 ) )   n = 50   d_n = 1 
assign Y[4'b1001] [51] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^51 ) )   n = 51   d_n = 1 
assign Y[4'b1001] [52] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^52 ) )   n = 52   d_n = 1 
assign Y[4'b1001] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^53 ) )   n = 53   d_n = 1 
assign Y[4'b1001] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^54 ) )   n = 54   d_n = 1 
assign Y[4'b1001] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^55 ) )   n = 55   d_n = 1 
assign Y[4'b1001] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^56 ) )   n = 56   d_n = 1 
assign Y[4'b1001] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^57 ) )   n = 57   d_n = 1 
assign Y[4'b1001] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^58 ) )   n = 58   d_n = 1 
assign Y[4'b1001] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^59 ) )   n = 59   d_n = 1 
assign Y[4'b1001] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^60 ) )   n = 60   d_n = 1 
assign Y[4'b1001] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^61 ) )   n = 61   d_n = 1 
assign Y[4'b1001] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^62 ) )   n = 62   d_n = 1 
assign Y[4'b1001] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^63 ) )   n = 63   d_n = 1 
assign Y[4'b1001] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  1 + 2^64 ) )   n = 64   d_n = 1 
assign Y[4'b1010] [01] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = -0 
assign Y[4'b1010] [02] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = -0 
assign Y[4'b1010] [03] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = -0 
assign Y[4'b1010] [04] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = -0 
assign Y[4'b1010] [05] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = -0 
assign Y[4'b1010] [06] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = -0 
assign Y[4'b1010] [07] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = -0 
assign Y[4'b1010] [08] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = -0 
assign Y[4'b1010] [09] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = -0 
assign Y[4'b1010] [10] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = -0 
assign Y[4'b1010] [11] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = -0 
assign Y[4'b1010] [12] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = -0 
assign Y[4'b1010] [13] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = -0 
assign Y[4'b1010] [14] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = -0 
assign Y[4'b1010] [15] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = -0 
assign Y[4'b1010] [16] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = -0 
assign Y[4'b1010] [17] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = -0 
assign Y[4'b1010] [18] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = -0 
assign Y[4'b1010] [19] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = -0 
assign Y[4'b1010] [20] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = -0 
assign Y[4'b1010] [21] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = -0 
assign Y[4'b1010] [22] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = -0 
assign Y[4'b1010] [23] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = -0 
assign Y[4'b1010] [24] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = -0 
assign Y[4'b1010] [25] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = -0 
assign Y[4'b1010] [26] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = -0 
assign Y[4'b1010] [27] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = -0 
assign Y[4'b1010] [28] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = -0 
assign Y[4'b1010] [29] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = -0 
assign Y[4'b1010] [30] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = -0 
assign Y[4'b1010] [31] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = -0 
assign Y[4'b1010] [32] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = -0 
assign Y[4'b1010] [33] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = -0 
assign Y[4'b1010] [34] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = -0 
assign Y[4'b1010] [35] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = -0 
assign Y[4'b1010] [36] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = -0 
assign Y[4'b1010] [37] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = -0 
assign Y[4'b1010] [38] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = -0 
assign Y[4'b1010] [39] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = -0 
assign Y[4'b1010] [40] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = -0 
assign Y[4'b1010] [41] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = -0 
assign Y[4'b1010] [42] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = -0 
assign Y[4'b1010] [43] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = -0 
assign Y[4'b1010] [44] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = -0 
assign Y[4'b1010] [45] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = -0 
assign Y[4'b1010] [46] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = -0 
assign Y[4'b1010] [47] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = -0 
assign Y[4'b1010] [48] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = -0 
assign Y[4'b1010] [49] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = -0 
assign Y[4'b1010] [50] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = -0 
assign Y[4'b1010] [51] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = -0 
assign Y[4'b1010] [52] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = -0 
assign Y[4'b1010] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = -0 
assign Y[4'b1010] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = -0 
assign Y[4'b1010] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = -0 
assign Y[4'b1010] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = -0 
assign Y[4'b1010] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = -0 
assign Y[4'b1010] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = -0 
assign Y[4'b1010] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = -0 
assign Y[4'b1010] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = -0 
assign Y[4'b1010] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = -0 
assign Y[4'b1010] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = -0 
assign Y[4'b1010] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = -0 
assign Y[4'b1010] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 +0.0000000000000000 =  0 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = -0 
assign Y[4'b1011] [01] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^1 ) )   n =  1   d_n = -1 
assign Y[4'b1011] [02] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^2 ) )   n =  2   d_n = -1 
assign Y[4'b1011] [03] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^3 ) )   n =  3   d_n = -1 
assign Y[4'b1011] [04] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^4 ) )   n =  4   d_n = -1 
assign Y[4'b1011] [05] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^5 ) )   n =  5   d_n = -1 
assign Y[4'b1011] [06] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^6 ) )   n =  6   d_n = -1 
assign Y[4'b1011] [07] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^7 ) )   n =  7   d_n = -1 
assign Y[4'b1011] [08] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^8 ) )   n =  8   d_n = -1 
assign Y[4'b1011] [09] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^9 ) )   n =  9   d_n = -1 
assign Y[4'b1011] [10] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^10 ) )   n = 10   d_n = -1 
assign Y[4'b1011] [11] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^11 ) )   n = 11   d_n = -1 
assign Y[4'b1011] [12] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^12 ) )   n = 12   d_n = -1 
assign Y[4'b1011] [13] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^13 ) )   n = 13   d_n = -1 
assign Y[4'b1011] [14] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^14 ) )   n = 14   d_n = -1 
assign Y[4'b1011] [15] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^15 ) )   n = 15   d_n = -1 
assign Y[4'b1011] [16] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^16 ) )   n = 16   d_n = -1 
assign Y[4'b1011] [17] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^17 ) )   n = 17   d_n = -1 
assign Y[4'b1011] [18] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^18 ) )   n = 18   d_n = -1 
assign Y[4'b1011] [19] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^19 ) )   n = 19   d_n = -1 
assign Y[4'b1011] [20] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^20 ) )   n = 20   d_n = -1 
assign Y[4'b1011] [21] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^21 ) )   n = 21   d_n = -1 
assign Y[4'b1011] [22] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^22 ) )   n = 22   d_n = -1 
assign Y[4'b1011] [23] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^23 ) )   n = 23   d_n = -1 
assign Y[4'b1011] [24] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^24 ) )   n = 24   d_n = -1 
assign Y[4'b1011] [25] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^25 ) )   n = 25   d_n = -1 
assign Y[4'b1011] [26] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^26 ) )   n = 26   d_n = -1 
assign Y[4'b1011] [27] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^27 ) )   n = 27   d_n = -1 
assign Y[4'b1011] [28] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^28 ) )   n = 28   d_n = -1 
assign Y[4'b1011] [29] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^29 ) )   n = 29   d_n = -1 
assign Y[4'b1011] [30] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^30 ) )   n = 30   d_n = -1 
assign Y[4'b1011] [31] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^31 ) )   n = 31   d_n = -1 
assign Y[4'b1011] [32] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^32 ) )   n = 32   d_n = -1 
assign Y[4'b1011] [33] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^33 ) )   n = 33   d_n = -1 
assign Y[4'b1011] [34] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^34 ) )   n = 34   d_n = -1 
assign Y[4'b1011] [35] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^35 ) )   n = 35   d_n = -1 
assign Y[4'b1011] [36] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^36 ) )   n = 36   d_n = -1 
assign Y[4'b1011] [37] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^37 ) )   n = 37   d_n = -1 
assign Y[4'b1011] [38] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^38 ) )   n = 38   d_n = -1 
assign Y[4'b1011] [39] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^39 ) )   n = 39   d_n = -1 
assign Y[4'b1011] [40] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^40 ) )   n = 40   d_n = -1 
assign Y[4'b1011] [41] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^41 ) )   n = 41   d_n = -1 
assign Y[4'b1011] [42] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^42 ) )   n = 42   d_n = -1 
assign Y[4'b1011] [43] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^43 ) )   n = 43   d_n = -1 
assign Y[4'b1011] [44] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^44 ) )   n = 44   d_n = -1 
assign Y[4'b1011] [45] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^45 ) )   n = 45   d_n = -1 
assign Y[4'b1011] [46] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^46 ) )   n = 46   d_n = -1 
assign Y[4'b1011] [47] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^47 ) )   n = 47   d_n = -1 
assign Y[4'b1011] [48] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^48 ) )   n = 48   d_n = -1 
assign Y[4'b1011] [49] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^49 ) )   n = 49   d_n = -1 
assign Y[4'b1011] [50] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^50 ) )   n = 50   d_n = -1 
assign Y[4'b1011] [51] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^51 ) )   n = 51   d_n = -1 
assign Y[4'b1011] [52] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^52 ) )   n = 52   d_n = -1 
assign Y[4'b1011] [53] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^53 ) )   n = 53   d_n = -1 
assign Y[4'b1011] [54] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^54 ) )   n = 54   d_n = -1 
assign Y[4'b1011] [55] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^55 ) )   n = 55   d_n = -1 
assign Y[4'b1011] [56] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^56 ) )   n = 56   d_n = -1 
assign Y[4'b1011] [57] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^57 ) )   n = 57   d_n = -1 
assign Y[4'b1011] [58] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^58 ) )   n = 58   d_n = -1 
assign Y[4'b1011] [59] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^59 ) )   n = 59   d_n = -1 
assign Y[4'b1011] [60] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^60 ) )   n = 60   d_n = -1 
assign Y[4'b1011] [61] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^61 ) )   n = 61   d_n = -1 
assign Y[4'b1011] [62] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^62 ) )   n = 62   d_n = -1 
assign Y[4'b1011] [63] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^63 ) )   n = 63   d_n = -1 
assign Y[4'b1011] [64] = 144'h 000000000000000000000000000000000000;  // 000000000000000000 -0.0000000000000000 =  0 * atan( 1 / ( -1 + 2^64 ) )   n = 64   d_n = -1 
assign Y[4'b1100] [01] = 144'h 000000201044421204021110204044880400;  // FFFC4A731F53C80000 -0.4636476090008061 = -1 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = -0-1i 
assign Y[4'b1100] [02] = 144'h 000000080044104044004221108002041000;  // FFFE0A48A06D380000 -0.2449786631268641 = -1 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = -0-1i 
assign Y[4'b1100] [03] = 144'h 000000020001110412220444440840104100;  // FFFF01522B2AA00000 -0.1243549945467614 = -1 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = -0-1i 
assign Y[4'b1100] [04] = 144'h 000000008000044441010412112000404880;  // FFFF802A9123500000 -0.0624188099959574 = -1 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = -0-1i 
assign Y[4'b1100] [05] = 144'h 000000002000001111104041222101102080;  // FFFFC0055488B00000 -0.0312398334302683 = -1 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = -0-1i 
assign Y[4'b1100] [06] = 144'h 000000000800000044444410101041088811;  // FFFFE000AAA4480000 -0.0156237286204768 = -1 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = -0-1i 
assign Y[4'b1100] [07] = 144'h 000000000200000001111111040404122210;  // FFFFF0001555200000 -0.0078123410601011 = -1 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = -0-1i 
assign Y[4'b1100] [08] = 144'h 000000000080000000044444444101010104;  // FFFFF80002AAA80000 -0.0039062301319670 = -1 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = -0-1i 
assign Y[4'b1100] [09] = 144'h 000000000020000000001111111110404040;  // FFFFFC000055580000 -0.0019531225164788 = -1 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = -0-1i 
assign Y[4'b1100] [10] = 144'h 000000000008000000000044444444441010;  // FFFFFE00000AA80000 -0.0009765621895593 = -1 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = -0-1i 
assign Y[4'b1100] [11] = 144'h 000000000002000000000001111111111104;  // FFFFFF000001580000 -0.0004882812111949 = -1 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = -0-1i 
assign Y[4'b1100] [12] = 144'h 000000000000800000000000044444444444;  // FFFFFF800000280000 -0.0002441406201494 = -1 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = -0-1i 
assign Y[4'b1100] [13] = 144'h 000000000000200000000000004888888888;  // FFFFFFC00000080000 -0.0001220703118937 = -1 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = -0-1i 
assign Y[4'b1100] [14] = 144'h 000000000000080000000000000122222222;  // FFFFFFE00000000000 -0.0000610351561742 = -1 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = -0-1i 
assign Y[4'b1100] [15] = 144'h 000000000000020000000000000004888888;  // FFFFFFF00000000000 -0.0000305175781155 = -1 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = -0-1i 
assign Y[4'b1100] [16] = 144'h 000000000000008000000000000000122222;  // FFFFFFF80000000000 -0.0000152587890613 = -1 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = -0-1i 
assign Y[4'b1100] [17] = 144'h 000000000000002000000000000000004888;  // FFFFFFFC0000000000 -0.0000076293945311 = -1 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = -0-1i 
assign Y[4'b1100] [18] = 144'h 000000000000000800000000000000000122;  // FFFFFFFE0000000000 -0.0000038146972656 = -1 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = -0-1i 
assign Y[4'b1100] [19] = 144'h 000000000000000200000000000000000004;  // FFFFFFFF0000000000 -0.0000019073486328 = -1 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = -0-1i 
assign Y[4'b1100] [20] = 144'h 000000000000000080000000000000000000;  // FFFFFFFF8000000000 -0.0000009536743164 = -1 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = -0-1i 
assign Y[4'b1100] [21] = 144'h 000000000000000020000000000000000000;  // FFFFFFFFC000000000 -0.0000004768371582 = -1 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = -0-1i 
assign Y[4'b1100] [22] = 144'h 000000000000000008000000000000000000;  // FFFFFFFFE000000000 -0.0000002384185791 = -1 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = -0-1i 
assign Y[4'b1100] [23] = 144'h 000000000000000002000000000000000000;  // FFFFFFFFF000000000 -0.0000001192092896 = -1 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = -0-1i 
assign Y[4'b1100] [24] = 144'h 000000000000000000800000000000000000;  // FFFFFFFFF800000000 -0.0000000596046448 = -1 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = -0-1i 
assign Y[4'b1100] [25] = 144'h 000000000000000000200000000000000000;  // FFFFFFFFFC00000000 -0.0000000298023224 = -1 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = -0-1i 
assign Y[4'b1100] [26] = 144'h 000000000000000000080000000000000000;  // FFFFFFFFFE00000000 -0.0000000149011612 = -1 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = -0-1i 
assign Y[4'b1100] [27] = 144'h 000000000000000000020000000000000000;  // FFFFFFFFFF00000000 -0.0000000074505806 = -1 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = -0-1i 
assign Y[4'b1100] [28] = 144'h 000000000000000000008000000000000000;  // FFFFFFFFFF80000000 -0.0000000037252903 = -1 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = -0-1i 
assign Y[4'b1100] [29] = 144'h 000000000000000000002000000000000000;  // FFFFFFFFFFC0000000 -0.0000000018626451 = -1 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = -0-1i 
assign Y[4'b1100] [30] = 144'h 000000000000000000000800000000000000;  // FFFFFFFFFFE0000000 -0.0000000009313226 = -1 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = -0-1i 
assign Y[4'b1100] [31] = 144'h 000000000000000000000200000000000000;  // FFFFFFFFFFF0000000 -0.0000000004656613 = -1 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = -0-1i 
assign Y[4'b1100] [32] = 144'h 000000000000000000000080000000000000;  // FFFFFFFFFFF8000000 -0.0000000002328306 = -1 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = -0-1i 
assign Y[4'b1100] [33] = 144'h 000000000000000000000020000000000000;  // FFFFFFFFFFFC000000 -0.0000000001164153 = -1 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = -0-1i 
assign Y[4'b1100] [34] = 144'h 000000000000000000000008000000000000;  // FFFFFFFFFFFE000000 -0.0000000000582077 = -1 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = -0-1i 
assign Y[4'b1100] [35] = 144'h 000000000000000000000002000000000000;  // FFFFFFFFFFFF000000 -0.0000000000291038 = -1 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = -0-1i 
assign Y[4'b1100] [36] = 144'h 000000000000000000000000800000000000;  // FFFFFFFFFFFF800000 -0.0000000000145519 = -1 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = -0-1i 
assign Y[4'b1100] [37] = 144'h 000000000000000000000000200000000000;  // FFFFFFFFFFFFC00000 -0.0000000000072760 = -1 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = -0-1i 
assign Y[4'b1100] [38] = 144'h 000000000000000000000000080000000000;  // FFFFFFFFFFFFE00000 -0.0000000000036380 = -1 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = -0-1i 
assign Y[4'b1100] [39] = 144'h 000000000000000000000000020000000000;  // FFFFFFFFFFFFF00000 -0.0000000000018190 = -1 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = -0-1i 
assign Y[4'b1100] [40] = 144'h 000000000000000000000000008000000000;  // FFFFFFFFFFFFF80000 -0.0000000000009095 = -1 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = -0-1i 
assign Y[4'b1100] [41] = 144'h 000000000000000000000000002000000000;  // 1000000000000000000 -0.0000000000004547 = -1 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = -0-1i 
assign Y[4'b1100] [42] = 144'h 000000000000000000000000000800000000;  // 1000000000000000000 -0.0000000000002274 = -1 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = -0-1i 
assign Y[4'b1100] [43] = 144'h 000000000000000000000000000200000000;  // 1000000000000000000 -0.0000000000001137 = -1 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = -0-1i 
assign Y[4'b1100] [44] = 144'h 000000000000000000000000000080000000;  // 1000000000000000000 -0.0000000000000568 = -1 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = -0-1i 
assign Y[4'b1100] [45] = 144'h 000000000000000000000000000020000000;  // 1000000000000000000 -0.0000000000000284 = -1 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = -0-1i 
assign Y[4'b1100] [46] = 144'h 000000000000000000000000000008000000;  // 1000000000000000000 -0.0000000000000142 = -1 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = -0-1i 
assign Y[4'b1100] [47] = 144'h 000000000000000000000000000002000000;  // 1000000000000000000 -0.0000000000000071 = -1 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = -0-1i 
assign Y[4'b1100] [48] = 144'h 000000000000000000000000000000800000;  // 1000000000000000000 -0.0000000000000036 = -1 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = -0-1i 
assign Y[4'b1100] [49] = 144'h 000000000000000000000000000000200000;  // 1000000000000000000 -0.0000000000000018 = -1 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = -0-1i 
assign Y[4'b1100] [50] = 144'h 000000000000000000000000000000080000;  // 1000000000000000000 -0.0000000000000009 = -1 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = -0-1i 
assign Y[4'b1100] [51] = 144'h 000000000000000000000000000000020000;  // 1000000000000000000 -0.0000000000000004 = -1 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = -0-1i 
assign Y[4'b1100] [52] = 144'h 000000000000000000000000000000008000;  // 1000000000000000000 -0.0000000000000002 = -1 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = -0-1i 
assign Y[4'b1100] [53] = 144'h 000000000000000000000000000000002000;  // 1000000000000000000 -0.0000000000000001 = -1 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = -0-1i 
assign Y[4'b1100] [54] = 144'h 000000000000000000000000000000000800;  // 1000000000000000000 -0.0000000000000001 = -1 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = -0-1i 
assign Y[4'b1100] [55] = 144'h 000000000000000000000000000000000200;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = -0-1i 
assign Y[4'b1100] [56] = 144'h 000000000000000000000000000000000080;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = -0-1i 
assign Y[4'b1100] [57] = 144'h 000000000000000000000000000000000020;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = -0-1i 
assign Y[4'b1100] [58] = 144'h 000000000000000000000000000000000008;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = -0-1i 
assign Y[4'b1100] [59] = 144'h 000000000000000000000000000000000002;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = -0-1i 
assign Y[4'b1100] [60] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = -0-1i 
assign Y[4'b1100] [61] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = -0-1i 
assign Y[4'b1100] [62] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = -0-1i 
assign Y[4'b1100] [63] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = -0-1i 
assign Y[4'b1100] [64] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = -0-1i 
assign Y[4'b1101] [01] = 144'h 000000088221010801208422122004100800;  // FFFD6D0E0B9B300000 -0.3217505543966422 = -1 * atan( 1 / (  1 + 2^1 ) )   n =  1   d_n = 1-1i 
assign Y[4'b1101] [02] = 144'h 000000084220202008004200410884021100;  // FFFE6BBBE070900000 -0.1973955598498807 = -1 * atan( 1 / (  1 + 2^2 ) )   n =  2   d_n = 1-1i 
assign Y[4'b1101] [03] = 144'h 000000020408880020021200020088084000;  // FFFF1D5FBF2FF00000 -0.1106572211738956 = -1 * atan( 1 / (  1 + 2^3 ) )   n =  3   d_n = 1-1i 
assign Y[4'b1101] [04] = 144'h 000000008040222200420080081004101200;  // FFFF87AB06F7E80000 -0.0587558227157227 = -1 * atan( 1 / (  1 + 2^4 ) )   n =  4   d_n = 1-1i 
assign Y[4'b1101] [05] = 144'h 000000002004008888804802000400104480;  // FFFFC1F5585F000000 -0.0302937599187751 = -1 * atan( 1 / (  1 + 2^5 ) )   n =  5   d_n = 1-1i 
assign Y[4'b1101] [06] = 144'h 000000000800400222222010842008044040;  // FFFFE07EAAC3980000 -0.0153834017805952 = -1 * atan( 1 / (  1 + 2^6 ) )   n =  6   d_n = 1-1i 
assign Y[4'b1101] [07] = 144'h 000000000200040008888888040080200044;  // FFFFF01FD556200000 -0.0077517827122069 = -1 * atan( 1 / (  1 + 2^7 ) )   n =  7   d_n = 1-1i 
assign Y[4'b1101] [08] = 144'h 000000000080004000222222220100484200;  // FFFFF807FAAAB00000 -0.0038910309466445 = -1 * atan( 1 / (  1 + 2^8 ) )   n =  8   d_n = 1-1i 
assign Y[4'b1101] [09] = 144'h 000000000020000400008888888880404808;  // FFFFFC01FF55580000 -0.0019493152697654 = -1 * atan( 1 / (  1 + 2^9 ) )   n =  9   d_n = 1-1i 
assign Y[4'b1101] [10] = 144'h 000000000008000040000222222222201010;  // FFFFFE007FEAA80000 -0.0009756094465646 = -1 * atan( 1 / (  1 + 2^10 ) )   n = 10   d_n = 1-1i 
assign Y[4'b1101] [11] = 144'h 000000000002000004000008888888888804;  // FFFFFF001FFD580000 -0.0004880429090311 = -1 * atan( 1 / (  1 + 2^11 ) )   n = 11   d_n = 1-1i 
assign Y[4'b1101] [12] = 144'h 000000000000800000400000222222222222;  // FFFFFF8007FFA80000 -0.0002440810300565 = -1 * atan( 1 / (  1 + 2^12 ) )   n = 12   d_n = 1-1i 
assign Y[4'b1101] [13] = 144'h 000000000000200000040000008888888888;  // FFFFFFC001FFF80000 -0.0001220554125515 = -1 * atan( 1 / (  1 + 2^13 ) )   n = 13   d_n = 1-1i 
assign Y[4'b1101] [14] = 144'h 000000000000080000004000000222222222;  // FFFFFFE00080000000 -0.0000610314311113 = -1 * atan( 1 / (  1 + 2^14 ) )   n = 14   d_n = 1-1i 
assign Y[4'b1101] [15] = 144'h 000000000000020000000400000008888888;  // FFFFFFF00020000000 -0.0000305166468214 = -1 * atan( 1 / (  1 + 2^15 ) )   n = 15   d_n = 1-1i 
assign Y[4'b1101] [16] = 144'h 000000000000008000000040000000222222;  // FFFFFFF80008000000 -0.0000152585562342 = -1 * atan( 1 / (  1 + 2^16 ) )   n = 16   d_n = 1-1i 
assign Y[4'b1101] [17] = 144'h 000000000000002000000004000000008888;  // FFFFFFFC0002000000 -0.0000076293363239 = -1 * atan( 1 / (  1 + 2^17 ) )   n = 17   d_n = 1-1i 
assign Y[4'b1101] [18] = 144'h 000000000000000800000000400000000222;  // FFFFFFFE0000800000 -0.0000038146827137 = -1 * atan( 1 / (  1 + 2^18 ) )   n = 18   d_n = 1-1i 
assign Y[4'b1101] [19] = 144'h 000000000000000200000000040000000008;  // FFFFFFFF0000200000 -0.0000019073449948 = -1 * atan( 1 / (  1 + 2^19 ) )   n = 19   d_n = 1-1i 
assign Y[4'b1101] [20] = 144'h 000000000000000080000000004000000000;  // FFFFFFFF8000080000 -0.0000009536734069 = -1 * atan( 1 / (  1 + 2^20 ) )   n = 20   d_n = 1-1i 
assign Y[4'b1101] [21] = 144'h 000000000000000020000000000400000000;  // FFFFFFFFC000000000 -0.0000004768369308 = -1 * atan( 1 / (  1 + 2^21 ) )   n = 21   d_n = 1-1i 
assign Y[4'b1101] [22] = 144'h 000000000000000008000000000040000000;  // FFFFFFFFE000000000 -0.0000002384185223 = -1 * atan( 1 / (  1 + 2^22 ) )   n = 22   d_n = 1-1i 
assign Y[4'b1101] [23] = 144'h 000000000000000002000000000004000000;  // FFFFFFFFF000000000 -0.0000001192092753 = -1 * atan( 1 / (  1 + 2^23 ) )   n = 23   d_n = 1-1i 
assign Y[4'b1101] [24] = 144'h 000000000000000000800000000000400000;  // FFFFFFFFF800000000 -0.0000000596046412 = -1 * atan( 1 / (  1 + 2^24 ) )   n = 24   d_n = 1-1i 
assign Y[4'b1101] [25] = 144'h 000000000000000000200000000000040000;  // FFFFFFFFFC00000000 -0.0000000298023215 = -1 * atan( 1 / (  1 + 2^25 ) )   n = 25   d_n = 1-1i 
assign Y[4'b1101] [26] = 144'h 000000000000000000080000000000004000;  // FFFFFFFFFE00000000 -0.0000000149011610 = -1 * atan( 1 / (  1 + 2^26 ) )   n = 26   d_n = 1-1i 
assign Y[4'b1101] [27] = 144'h 000000000000000000020000000000000400;  // FFFFFFFFFF00000000 -0.0000000074505805 = -1 * atan( 1 / (  1 + 2^27 ) )   n = 27   d_n = 1-1i 
assign Y[4'b1101] [28] = 144'h 000000000000000000008000000000000040;  // FFFFFFFFFF80000000 -0.0000000037252903 = -1 * atan( 1 / (  1 + 2^28 ) )   n = 28   d_n = 1-1i 
assign Y[4'b1101] [29] = 144'h 000000000000000000002000000000000004;  // FFFFFFFFFFC0000000 -0.0000000018626451 = -1 * atan( 1 / (  1 + 2^29 ) )   n = 29   d_n = 1-1i 
assign Y[4'b1101] [30] = 144'h 000000000000000000000800000000000000;  // FFFFFFFFFFE0000000 -0.0000000009313226 = -1 * atan( 1 / (  1 + 2^30 ) )   n = 30   d_n = 1-1i 
assign Y[4'b1101] [31] = 144'h 000000000000000000000200000000000000;  // FFFFFFFFFFF0000000 -0.0000000004656613 = -1 * atan( 1 / (  1 + 2^31 ) )   n = 31   d_n = 1-1i 
assign Y[4'b1101] [32] = 144'h 000000000000000000000080000000000000;  // FFFFFFFFFFF8000000 -0.0000000002328306 = -1 * atan( 1 / (  1 + 2^32 ) )   n = 32   d_n = 1-1i 
assign Y[4'b1101] [33] = 144'h 000000000000000000000020000000000000;  // FFFFFFFFFFFC000000 -0.0000000001164153 = -1 * atan( 1 / (  1 + 2^33 ) )   n = 33   d_n = 1-1i 
assign Y[4'b1101] [34] = 144'h 000000000000000000000008000000000000;  // FFFFFFFFFFFE000000 -0.0000000000582077 = -1 * atan( 1 / (  1 + 2^34 ) )   n = 34   d_n = 1-1i 
assign Y[4'b1101] [35] = 144'h 000000000000000000000002000000000000;  // FFFFFFFFFFFF000000 -0.0000000000291038 = -1 * atan( 1 / (  1 + 2^35 ) )   n = 35   d_n = 1-1i 
assign Y[4'b1101] [36] = 144'h 000000000000000000000000800000000000;  // FFFFFFFFFFFF800000 -0.0000000000145519 = -1 * atan( 1 / (  1 + 2^36 ) )   n = 36   d_n = 1-1i 
assign Y[4'b1101] [37] = 144'h 000000000000000000000000200000000000;  // FFFFFFFFFFFFC00000 -0.0000000000072760 = -1 * atan( 1 / (  1 + 2^37 ) )   n = 37   d_n = 1-1i 
assign Y[4'b1101] [38] = 144'h 000000000000000000000000080000000000;  // FFFFFFFFFFFFE00000 -0.0000000000036380 = -1 * atan( 1 / (  1 + 2^38 ) )   n = 38   d_n = 1-1i 
assign Y[4'b1101] [39] = 144'h 000000000000000000000000020000000000;  // FFFFFFFFFFFFF00000 -0.0000000000018190 = -1 * atan( 1 / (  1 + 2^39 ) )   n = 39   d_n = 1-1i 
assign Y[4'b1101] [40] = 144'h 000000000000000000000000008000000000;  // FFFFFFFFFFFFF80000 -0.0000000000009095 = -1 * atan( 1 / (  1 + 2^40 ) )   n = 40   d_n = 1-1i 
assign Y[4'b1101] [41] = 144'h 000000000000000000000000002000000000;  // 1000000000000000000 -0.0000000000004547 = -1 * atan( 1 / (  1 + 2^41 ) )   n = 41   d_n = 1-1i 
assign Y[4'b1101] [42] = 144'h 000000000000000000000000000800000000;  // 1000000000000000000 -0.0000000000002274 = -1 * atan( 1 / (  1 + 2^42 ) )   n = 42   d_n = 1-1i 
assign Y[4'b1101] [43] = 144'h 000000000000000000000000000200000000;  // 1000000000000000000 -0.0000000000001137 = -1 * atan( 1 / (  1 + 2^43 ) )   n = 43   d_n = 1-1i 
assign Y[4'b1101] [44] = 144'h 000000000000000000000000000080000000;  // 1000000000000000000 -0.0000000000000568 = -1 * atan( 1 / (  1 + 2^44 ) )   n = 44   d_n = 1-1i 
assign Y[4'b1101] [45] = 144'h 000000000000000000000000000020000000;  // 1000000000000000000 -0.0000000000000284 = -1 * atan( 1 / (  1 + 2^45 ) )   n = 45   d_n = 1-1i 
assign Y[4'b1101] [46] = 144'h 000000000000000000000000000008000000;  // 1000000000000000000 -0.0000000000000142 = -1 * atan( 1 / (  1 + 2^46 ) )   n = 46   d_n = 1-1i 
assign Y[4'b1101] [47] = 144'h 000000000000000000000000000002000000;  // 1000000000000000000 -0.0000000000000071 = -1 * atan( 1 / (  1 + 2^47 ) )   n = 47   d_n = 1-1i 
assign Y[4'b1101] [48] = 144'h 000000000000000000000000000000800000;  // 1000000000000000000 -0.0000000000000036 = -1 * atan( 1 / (  1 + 2^48 ) )   n = 48   d_n = 1-1i 
assign Y[4'b1101] [49] = 144'h 000000000000000000000000000000200000;  // 1000000000000000000 -0.0000000000000018 = -1 * atan( 1 / (  1 + 2^49 ) )   n = 49   d_n = 1-1i 
assign Y[4'b1101] [50] = 144'h 000000000000000000000000000000080000;  // 1000000000000000000 -0.0000000000000009 = -1 * atan( 1 / (  1 + 2^50 ) )   n = 50   d_n = 1-1i 
assign Y[4'b1101] [51] = 144'h 000000000000000000000000000000020000;  // 1000000000000000000 -0.0000000000000004 = -1 * atan( 1 / (  1 + 2^51 ) )   n = 51   d_n = 1-1i 
assign Y[4'b1101] [52] = 144'h 000000000000000000000000000000008000;  // 1000000000000000000 -0.0000000000000002 = -1 * atan( 1 / (  1 + 2^52 ) )   n = 52   d_n = 1-1i 
assign Y[4'b1101] [53] = 144'h 000000000000000000000000000000002000;  // 1000000000000000000 -0.0000000000000001 = -1 * atan( 1 / (  1 + 2^53 ) )   n = 53   d_n = 1-1i 
assign Y[4'b1101] [54] = 144'h 000000000000000000000000000000000800;  // 1000000000000000000 -0.0000000000000001 = -1 * atan( 1 / (  1 + 2^54 ) )   n = 54   d_n = 1-1i 
assign Y[4'b1101] [55] = 144'h 000000000000000000000000000000000200;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^55 ) )   n = 55   d_n = 1-1i 
assign Y[4'b1101] [56] = 144'h 000000000000000000000000000000000080;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^56 ) )   n = 56   d_n = 1-1i 
assign Y[4'b1101] [57] = 144'h 000000000000000000000000000000000020;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^57 ) )   n = 57   d_n = 1-1i 
assign Y[4'b1101] [58] = 144'h 000000000000000000000000000000000008;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^58 ) )   n = 58   d_n = 1-1i 
assign Y[4'b1101] [59] = 144'h 000000000000000000000000000000000002;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^59 ) )   n = 59   d_n = 1-1i 
assign Y[4'b1101] [60] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^60 ) )   n = 60   d_n = 1-1i 
assign Y[4'b1101] [61] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^61 ) )   n = 61   d_n = 1-1i 
assign Y[4'b1101] [62] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^62 ) )   n = 62   d_n = 1-1i 
assign Y[4'b1101] [63] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^63 ) )   n = 63   d_n = 1-1i 
assign Y[4'b1101] [64] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  1 + 2^64 ) )   n = 64   d_n = 1-1i 
assign Y[4'b1110] [01] = 144'h 000000201044421204021110204044880400;  // FFFC4A731F53C80000 -0.4636476090008061 = -1 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = -0-1i 
assign Y[4'b1110] [02] = 144'h 000000080044104044004221108002041000;  // FFFE0A48A06D380000 -0.2449786631268641 = -1 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = -0-1i 
assign Y[4'b1110] [03] = 144'h 000000020001110412220444440840104100;  // FFFF01522B2AA00000 -0.1243549945467614 = -1 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = -0-1i 
assign Y[4'b1110] [04] = 144'h 000000008000044441010412112000404880;  // FFFF802A9123500000 -0.0624188099959574 = -1 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = -0-1i 
assign Y[4'b1110] [05] = 144'h 000000002000001111104041222101102080;  // FFFFC0055488B00000 -0.0312398334302683 = -1 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = -0-1i 
assign Y[4'b1110] [06] = 144'h 000000000800000044444410101041088811;  // FFFFE000AAA4480000 -0.0156237286204768 = -1 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = -0-1i 
assign Y[4'b1110] [07] = 144'h 000000000200000001111111040404122210;  // FFFFF0001555200000 -0.0078123410601011 = -1 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = -0-1i 
assign Y[4'b1110] [08] = 144'h 000000000080000000044444444101010104;  // FFFFF80002AAA80000 -0.0039062301319670 = -1 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = -0-1i 
assign Y[4'b1110] [09] = 144'h 000000000020000000001111111110404040;  // FFFFFC000055580000 -0.0019531225164788 = -1 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = -0-1i 
assign Y[4'b1110] [10] = 144'h 000000000008000000000044444444441010;  // FFFFFE00000AA80000 -0.0009765621895593 = -1 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = -0-1i 
assign Y[4'b1110] [11] = 144'h 000000000002000000000001111111111104;  // FFFFFF000001580000 -0.0004882812111949 = -1 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = -0-1i 
assign Y[4'b1110] [12] = 144'h 000000000000800000000000044444444444;  // FFFFFF800000280000 -0.0002441406201494 = -1 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = -0-1i 
assign Y[4'b1110] [13] = 144'h 000000000000200000000000004888888888;  // FFFFFFC00000080000 -0.0001220703118937 = -1 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = -0-1i 
assign Y[4'b1110] [14] = 144'h 000000000000080000000000000122222222;  // FFFFFFE00000000000 -0.0000610351561742 = -1 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = -0-1i 
assign Y[4'b1110] [15] = 144'h 000000000000020000000000000004888888;  // FFFFFFF00000000000 -0.0000305175781155 = -1 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = -0-1i 
assign Y[4'b1110] [16] = 144'h 000000000000008000000000000000122222;  // FFFFFFF80000000000 -0.0000152587890613 = -1 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = -0-1i 
assign Y[4'b1110] [17] = 144'h 000000000000002000000000000000004888;  // FFFFFFFC0000000000 -0.0000076293945311 = -1 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = -0-1i 
assign Y[4'b1110] [18] = 144'h 000000000000000800000000000000000122;  // FFFFFFFE0000000000 -0.0000038146972656 = -1 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = -0-1i 
assign Y[4'b1110] [19] = 144'h 000000000000000200000000000000000004;  // FFFFFFFF0000000000 -0.0000019073486328 = -1 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = -0-1i 
assign Y[4'b1110] [20] = 144'h 000000000000000080000000000000000000;  // FFFFFFFF8000000000 -0.0000009536743164 = -1 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = -0-1i 
assign Y[4'b1110] [21] = 144'h 000000000000000020000000000000000000;  // FFFFFFFFC000000000 -0.0000004768371582 = -1 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = -0-1i 
assign Y[4'b1110] [22] = 144'h 000000000000000008000000000000000000;  // FFFFFFFFE000000000 -0.0000002384185791 = -1 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = -0-1i 
assign Y[4'b1110] [23] = 144'h 000000000000000002000000000000000000;  // FFFFFFFFF000000000 -0.0000001192092896 = -1 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = -0-1i 
assign Y[4'b1110] [24] = 144'h 000000000000000000800000000000000000;  // FFFFFFFFF800000000 -0.0000000596046448 = -1 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = -0-1i 
assign Y[4'b1110] [25] = 144'h 000000000000000000200000000000000000;  // FFFFFFFFFC00000000 -0.0000000298023224 = -1 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = -0-1i 
assign Y[4'b1110] [26] = 144'h 000000000000000000080000000000000000;  // FFFFFFFFFE00000000 -0.0000000149011612 = -1 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = -0-1i 
assign Y[4'b1110] [27] = 144'h 000000000000000000020000000000000000;  // FFFFFFFFFF00000000 -0.0000000074505806 = -1 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = -0-1i 
assign Y[4'b1110] [28] = 144'h 000000000000000000008000000000000000;  // FFFFFFFFFF80000000 -0.0000000037252903 = -1 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = -0-1i 
assign Y[4'b1110] [29] = 144'h 000000000000000000002000000000000000;  // FFFFFFFFFFC0000000 -0.0000000018626451 = -1 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = -0-1i 
assign Y[4'b1110] [30] = 144'h 000000000000000000000800000000000000;  // FFFFFFFFFFE0000000 -0.0000000009313226 = -1 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = -0-1i 
assign Y[4'b1110] [31] = 144'h 000000000000000000000200000000000000;  // FFFFFFFFFFF0000000 -0.0000000004656613 = -1 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = -0-1i 
assign Y[4'b1110] [32] = 144'h 000000000000000000000080000000000000;  // FFFFFFFFFFF8000000 -0.0000000002328306 = -1 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = -0-1i 
assign Y[4'b1110] [33] = 144'h 000000000000000000000020000000000000;  // FFFFFFFFFFFC000000 -0.0000000001164153 = -1 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = -0-1i 
assign Y[4'b1110] [34] = 144'h 000000000000000000000008000000000000;  // FFFFFFFFFFFE000000 -0.0000000000582077 = -1 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = -0-1i 
assign Y[4'b1110] [35] = 144'h 000000000000000000000002000000000000;  // FFFFFFFFFFFF000000 -0.0000000000291038 = -1 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = -0-1i 
assign Y[4'b1110] [36] = 144'h 000000000000000000000000800000000000;  // FFFFFFFFFFFF800000 -0.0000000000145519 = -1 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = -0-1i 
assign Y[4'b1110] [37] = 144'h 000000000000000000000000200000000000;  // FFFFFFFFFFFFC00000 -0.0000000000072760 = -1 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = -0-1i 
assign Y[4'b1110] [38] = 144'h 000000000000000000000000080000000000;  // FFFFFFFFFFFFE00000 -0.0000000000036380 = -1 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = -0-1i 
assign Y[4'b1110] [39] = 144'h 000000000000000000000000020000000000;  // FFFFFFFFFFFFF00000 -0.0000000000018190 = -1 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = -0-1i 
assign Y[4'b1110] [40] = 144'h 000000000000000000000000008000000000;  // FFFFFFFFFFFFF80000 -0.0000000000009095 = -1 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = -0-1i 
assign Y[4'b1110] [41] = 144'h 000000000000000000000000002000000000;  // 1000000000000000000 -0.0000000000004547 = -1 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = -0-1i 
assign Y[4'b1110] [42] = 144'h 000000000000000000000000000800000000;  // 1000000000000000000 -0.0000000000002274 = -1 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = -0-1i 
assign Y[4'b1110] [43] = 144'h 000000000000000000000000000200000000;  // 1000000000000000000 -0.0000000000001137 = -1 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = -0-1i 
assign Y[4'b1110] [44] = 144'h 000000000000000000000000000080000000;  // 1000000000000000000 -0.0000000000000568 = -1 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = -0-1i 
assign Y[4'b1110] [45] = 144'h 000000000000000000000000000020000000;  // 1000000000000000000 -0.0000000000000284 = -1 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = -0-1i 
assign Y[4'b1110] [46] = 144'h 000000000000000000000000000008000000;  // 1000000000000000000 -0.0000000000000142 = -1 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = -0-1i 
assign Y[4'b1110] [47] = 144'h 000000000000000000000000000002000000;  // 1000000000000000000 -0.0000000000000071 = -1 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = -0-1i 
assign Y[4'b1110] [48] = 144'h 000000000000000000000000000000800000;  // 1000000000000000000 -0.0000000000000036 = -1 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = -0-1i 
assign Y[4'b1110] [49] = 144'h 000000000000000000000000000000200000;  // 1000000000000000000 -0.0000000000000018 = -1 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = -0-1i 
assign Y[4'b1110] [50] = 144'h 000000000000000000000000000000080000;  // 1000000000000000000 -0.0000000000000009 = -1 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = -0-1i 
assign Y[4'b1110] [51] = 144'h 000000000000000000000000000000020000;  // 1000000000000000000 -0.0000000000000004 = -1 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = -0-1i 
assign Y[4'b1110] [52] = 144'h 000000000000000000000000000000008000;  // 1000000000000000000 -0.0000000000000002 = -1 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = -0-1i 
assign Y[4'b1110] [53] = 144'h 000000000000000000000000000000002000;  // 1000000000000000000 -0.0000000000000001 = -1 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = -0-1i 
assign Y[4'b1110] [54] = 144'h 000000000000000000000000000000000800;  // 1000000000000000000 -0.0000000000000001 = -1 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = -0-1i 
assign Y[4'b1110] [55] = 144'h 000000000000000000000000000000000200;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = -0-1i 
assign Y[4'b1110] [56] = 144'h 000000000000000000000000000000000080;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = -0-1i 
assign Y[4'b1110] [57] = 144'h 000000000000000000000000000000000020;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = -0-1i 
assign Y[4'b1110] [58] = 144'h 000000000000000000000000000000000008;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = -0-1i 
assign Y[4'b1110] [59] = 144'h 000000000000000000000000000000000002;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = -0-1i 
assign Y[4'b1110] [60] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = -0-1i 
assign Y[4'b1110] [61] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = -0-1i 
assign Y[4'b1110] [62] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = -0-1i 
assign Y[4'b1110] [63] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = -0-1i 
assign Y[4'b1110] [64] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = -0-1i 
assign Y[4'b1111] [01] = 144'h 000000842080800112220202021120840000;  // FFF9B7812AEEF80000 -0.7853981633974483 = -1 * atan( 1 / ( -1 + 2^1 ) )   n =  1   d_n = -1-1i 
assign Y[4'b1111] [02] = 144'h 000000088221010801208422122004100800;  // FFFD6D0E0B9B300000 -0.3217505543966422 = -1 * atan( 1 / ( -1 + 2^2 ) )   n =  2   d_n = -1-1i 
assign Y[4'b1111] [03] = 144'h 000000020808881101102080442042041200;  // FFFEDD6513B8A00000 -0.1418970546041639 = -1 * atan( 1 / ( -1 + 2^3 ) )   n =  3   d_n = -1-1i 
assign Y[4'b1111] [04] = 144'h 000000008080222204201121004810420800;  // FFFF77AB1C4D080000 -0.0665681637758238 = -1 * atan( 1 / ( -1 + 2^4 ) )   n =  4   d_n = -1-1i 
assign Y[4'b1111] [05] = 144'h 000000002008008888812210488211210400;  // FFFFBDF558B4580000 -0.0322468824352539 = -1 * atan( 1 / ( -1 + 2^5 ) )   n =  5   d_n = -1-1i 
assign Y[4'b1111] [06] = 144'h 000000000800800222222011020110800880;  // FFFFDF7EAAC4F00000 -0.0158716829917901 = -1 * atan( 1 / ( -1 + 2^6 ) )   n =  6   d_n = -1-1i 
assign Y[4'b1111] [07] = 144'h 000000000200080008888888041121048802;  // FFFFEFDFD556280000 -0.0078738530241005 = -1 * atan( 1 / ( -1 + 2^7 ) )   n =  7   d_n = -1-1i 
assign Y[4'b1111] [08] = 144'h 000000000080008000222222220104202011;  // FFFFF7F7FAAAB00000 -0.0039215485247600 = -1 * atan( 1 / ( -1 + 2^8 ) )   n =  8   d_n = -1-1i 
assign Y[4'b1111] [09] = 144'h 000000000020000800008888888880412212;  // FFFFFBFDFF55580000 -0.0019569446642965 = -1 * atan( 1 / ( -1 + 2^9 ) )   n =  9   d_n = -1-1i 
assign Y[4'b1111] [10] = 144'h 000000000008000080000222222222201011;  // FFFFFDFF7FEAA80000 -0.0009775167951974 = -1 * atan( 1 / ( -1 + 2^10 ) )   n = 10   d_n = -1-1i 
assign Y[4'b1111] [11] = 144'h 000000000002000008000008888888888804;  // FFFFFEFFDFFD580000 -0.0004885197461893 = -1 * atan( 1 / ( -1 + 2^11 ) )   n = 11   d_n = -1-1i 
assign Y[4'b1111] [12] = 144'h 000000000000800000800000222222222222;  // FFFFFF7FF7FFA80000 -0.0002442002393461 = -1 * atan( 1 / ( -1 + 2^12 ) )   n = 12   d_n = -1-1i 
assign Y[4'b1111] [13] = 144'h 000000000000200000080000008888888888;  // FFFFFFBFFDFFF80000 -0.0001220852148739 = -1 * atan( 1 / ( -1 + 2^13 ) )   n = 13   d_n = -1-1i 
assign Y[4'b1111] [14] = 144'h 000000000000080000008000000222222222;  // FFFFFFDFFF80000000 -0.0000610388816919 = -1 * atan( 1 / ( -1 + 2^14 ) )   n = 14   d_n = -1-1i 
assign Y[4'b1111] [15] = 144'h 000000000000020000000800000008888888;  // FFFFFFEFFFE0000000 -0.0000305185094665 = -1 * atan( 1 / ( -1 + 2^15 ) )   n = 15   d_n = -1-1i 
assign Y[4'b1111] [16] = 144'h 000000000000008000000080000000222222;  // FFFFFFF7FFF8000000 -0.0000152590218955 = -1 * atan( 1 / ( -1 + 2^16 ) )   n = 16   d_n = -1-1i 
assign Y[4'b1111] [17] = 144'h 000000000000002000000008000000008888;  // FFFFFFFBFFFE000000 -0.0000076294527392 = -1 * atan( 1 / ( -1 + 2^17 ) )   n = 17   d_n = -1-1i 
assign Y[4'b1111] [18] = 144'h 000000000000000800000000800000000222;  // FFFFFFFDFFFF800000 -0.0000038147118176 = -1 * atan( 1 / ( -1 + 2^18 ) )   n = 18   d_n = -1-1i 
assign Y[4'b1111] [19] = 144'h 000000000000000200000000080000000008;  // FFFFFFFEFFFFE00000 -0.0000019073522708 = -1 * atan( 1 / ( -1 + 2^19 ) )   n = 19   d_n = -1-1i 
assign Y[4'b1111] [20] = 144'h 000000000000000080000000008000000000;  // FFFFFFFF7FFFF80000 -0.0000009536752259 = -1 * atan( 1 / ( -1 + 2^20 ) )   n = 20   d_n = -1-1i 
assign Y[4'b1111] [21] = 144'h 000000000000000020000000000800000000;  // FFFFFFFFC000000000 -0.0000004768373856 = -1 * atan( 1 / ( -1 + 2^21 ) )   n = 21   d_n = -1-1i 
assign Y[4'b1111] [22] = 144'h 000000000000000008000000000080000000;  // FFFFFFFFE000000000 -0.0000002384186359 = -1 * atan( 1 / ( -1 + 2^22 ) )   n = 22   d_n = -1-1i 
assign Y[4'b1111] [23] = 144'h 000000000000000002000000000008000000;  // FFFFFFFFF000000000 -0.0000001192093038 = -1 * atan( 1 / ( -1 + 2^23 ) )   n = 23   d_n = -1-1i 
assign Y[4'b1111] [24] = 144'h 000000000000000000800000000000800000;  // FFFFFFFFF800000000 -0.0000000596046483 = -1 * atan( 1 / ( -1 + 2^24 ) )   n = 24   d_n = -1-1i 
assign Y[4'b1111] [25] = 144'h 000000000000000000200000000000080000;  // FFFFFFFFFC00000000 -0.0000000298023233 = -1 * atan( 1 / ( -1 + 2^25 ) )   n = 25   d_n = -1-1i 
assign Y[4'b1111] [26] = 144'h 000000000000000000080000000000008000;  // FFFFFFFFFE00000000 -0.0000000149011614 = -1 * atan( 1 / ( -1 + 2^26 ) )   n = 26   d_n = -1-1i 
assign Y[4'b1111] [27] = 144'h 000000000000000000020000000000000800;  // FFFFFFFFFF00000000 -0.0000000074505807 = -1 * atan( 1 / ( -1 + 2^27 ) )   n = 27   d_n = -1-1i 
assign Y[4'b1111] [28] = 144'h 000000000000000000008000000000000080;  // FFFFFFFFFF80000000 -0.0000000037252903 = -1 * atan( 1 / ( -1 + 2^28 ) )   n = 28   d_n = -1-1i 
assign Y[4'b1111] [29] = 144'h 000000000000000000002000000000000008;  // FFFFFFFFFFC0000000 -0.0000000018626452 = -1 * atan( 1 / ( -1 + 2^29 ) )   n = 29   d_n = -1-1i 
assign Y[4'b1111] [30] = 144'h 000000000000000000000800000000000000;  // FFFFFFFFFFE0000000 -0.0000000009313226 = -1 * atan( 1 / ( -1 + 2^30 ) )   n = 30   d_n = -1-1i 
assign Y[4'b1111] [31] = 144'h 000000000000000000000200000000000000;  // FFFFFFFFFFF0000000 -0.0000000004656613 = -1 * atan( 1 / ( -1 + 2^31 ) )   n = 31   d_n = -1-1i 
assign Y[4'b1111] [32] = 144'h 000000000000000000000080000000000000;  // FFFFFFFFFFF8000000 -0.0000000002328306 = -1 * atan( 1 / ( -1 + 2^32 ) )   n = 32   d_n = -1-1i 
assign Y[4'b1111] [33] = 144'h 000000000000000000000020000000000000;  // FFFFFFFFFFFC000000 -0.0000000001164153 = -1 * atan( 1 / ( -1 + 2^33 ) )   n = 33   d_n = -1-1i 
assign Y[4'b1111] [34] = 144'h 000000000000000000000008000000000000;  // FFFFFFFFFFFE000000 -0.0000000000582077 = -1 * atan( 1 / ( -1 + 2^34 ) )   n = 34   d_n = -1-1i 
assign Y[4'b1111] [35] = 144'h 000000000000000000000002000000000000;  // FFFFFFFFFFFF000000 -0.0000000000291038 = -1 * atan( 1 / ( -1 + 2^35 ) )   n = 35   d_n = -1-1i 
assign Y[4'b1111] [36] = 144'h 000000000000000000000000800000000000;  // FFFFFFFFFFFF800000 -0.0000000000145519 = -1 * atan( 1 / ( -1 + 2^36 ) )   n = 36   d_n = -1-1i 
assign Y[4'b1111] [37] = 144'h 000000000000000000000000200000000000;  // FFFFFFFFFFFFC00000 -0.0000000000072760 = -1 * atan( 1 / ( -1 + 2^37 ) )   n = 37   d_n = -1-1i 
assign Y[4'b1111] [38] = 144'h 000000000000000000000000080000000000;  // FFFFFFFFFFFFE00000 -0.0000000000036380 = -1 * atan( 1 / ( -1 + 2^38 ) )   n = 38   d_n = -1-1i 
assign Y[4'b1111] [39] = 144'h 000000000000000000000000020000000000;  // FFFFFFFFFFFFF00000 -0.0000000000018190 = -1 * atan( 1 / ( -1 + 2^39 ) )   n = 39   d_n = -1-1i 
assign Y[4'b1111] [40] = 144'h 000000000000000000000000008000000000;  // FFFFFFFFFFFFF80000 -0.0000000000009095 = -1 * atan( 1 / ( -1 + 2^40 ) )   n = 40   d_n = -1-1i 
assign Y[4'b1111] [41] = 144'h 000000000000000000000000002000000000;  // FFFFFFFFFFFFF80000 -0.0000000000004547 = -1 * atan( 1 / ( -1 + 2^41 ) )   n = 41   d_n = -1-1i 
assign Y[4'b1111] [42] = 144'h 000000000000000000000000000800000000;  // 1000000000000000000 -0.0000000000002274 = -1 * atan( 1 / ( -1 + 2^42 ) )   n = 42   d_n = -1-1i 
assign Y[4'b1111] [43] = 144'h 000000000000000000000000000200000000;  // 1000000000000000000 -0.0000000000001137 = -1 * atan( 1 / ( -1 + 2^43 ) )   n = 43   d_n = -1-1i 
assign Y[4'b1111] [44] = 144'h 000000000000000000000000000080000000;  // 1000000000000000000 -0.0000000000000568 = -1 * atan( 1 / ( -1 + 2^44 ) )   n = 44   d_n = -1-1i 
assign Y[4'b1111] [45] = 144'h 000000000000000000000000000020000000;  // 1000000000000000000 -0.0000000000000284 = -1 * atan( 1 / ( -1 + 2^45 ) )   n = 45   d_n = -1-1i 
assign Y[4'b1111] [46] = 144'h 000000000000000000000000000008000000;  // 1000000000000000000 -0.0000000000000142 = -1 * atan( 1 / ( -1 + 2^46 ) )   n = 46   d_n = -1-1i 
assign Y[4'b1111] [47] = 144'h 000000000000000000000000000002000000;  // 1000000000000000000 -0.0000000000000071 = -1 * atan( 1 / ( -1 + 2^47 ) )   n = 47   d_n = -1-1i 
assign Y[4'b1111] [48] = 144'h 000000000000000000000000000000800000;  // 1000000000000000000 -0.0000000000000036 = -1 * atan( 1 / ( -1 + 2^48 ) )   n = 48   d_n = -1-1i 
assign Y[4'b1111] [49] = 144'h 000000000000000000000000000000200000;  // 1000000000000000000 -0.0000000000000018 = -1 * atan( 1 / ( -1 + 2^49 ) )   n = 49   d_n = -1-1i 
assign Y[4'b1111] [50] = 144'h 000000000000000000000000000000080000;  // 1000000000000000000 -0.0000000000000009 = -1 * atan( 1 / ( -1 + 2^50 ) )   n = 50   d_n = -1-1i 
assign Y[4'b1111] [51] = 144'h 000000000000000000000000000000020000;  // 1000000000000000000 -0.0000000000000004 = -1 * atan( 1 / ( -1 + 2^51 ) )   n = 51   d_n = -1-1i 
assign Y[4'b1111] [52] = 144'h 000000000000000000000000000000008000;  // 1000000000000000000 -0.0000000000000002 = -1 * atan( 1 / ( -1 + 2^52 ) )   n = 52   d_n = -1-1i 
assign Y[4'b1111] [53] = 144'h 000000000000000000000000000000002000;  // 1000000000000000000 -0.0000000000000001 = -1 * atan( 1 / ( -1 + 2^53 ) )   n = 53   d_n = -1-1i 
assign Y[4'b1111] [54] = 144'h 000000000000000000000000000000000800;  // 1000000000000000000 -0.0000000000000001 = -1 * atan( 1 / ( -1 + 2^54 ) )   n = 54   d_n = -1-1i 
assign Y[4'b1111] [55] = 144'h 000000000000000000000000000000000200;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^55 ) )   n = 55   d_n = -1-1i 
assign Y[4'b1111] [56] = 144'h 000000000000000000000000000000000080;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^56 ) )   n = 56   d_n = -1-1i 
assign Y[4'b1111] [57] = 144'h 000000000000000000000000000000000020;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^57 ) )   n = 57   d_n = -1-1i 
assign Y[4'b1111] [58] = 144'h 000000000000000000000000000000000008;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^58 ) )   n = 58   d_n = -1-1i 
assign Y[4'b1111] [59] = 144'h 000000000000000000000000000000000002;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^59 ) )   n = 59   d_n = -1-1i 
assign Y[4'b1111] [60] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^60 ) )   n = 60   d_n = -1-1i 
assign Y[4'b1111] [61] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^61 ) )   n = 61   d_n = -1-1i 
assign Y[4'b1111] [62] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^62 ) )   n = 62   d_n = -1-1i 
assign Y[4'b1111] [63] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^63 ) )   n = 63   d_n = -1-1i 
assign Y[4'b1111] [64] = 144'h 000000000000000000000000000000000000;  // 1000000000000000000 -0.0000000000000000 = -1 * atan( 1 / ( -1 + 2^64 ) )   n = 64   d_n = -1-1i 
//
//
//--------------------------------------------------------------------------------
// This LUT uses 22 bits which represent 22 twos complement digits. 
// They are represented by 6 hexadecimal digits. 
// After the LUT value you have the floating point representation. 
// Since we use 14 bits for the integer part then the first 4.0 hexa digits represent the integer part. 
// The rest 2.0 hexa digits represent the fractional part.
// Example:
//sign u[4'bXXXX] [XX] = 22'h 000000;  //   +0.0000000000000001
//--------------------------------------------------------------------------------
//
assign u[4'b0000] [01] = 22'h 000000;  // +0.0000000000000000 = 2^ 1 * ln( 1 +  0 * 2^(- 1+1) + ( 0^2+ 0^2) * 2^(-2* 1) )   n =  1   d_n = 0 
assign u[4'b0000] [02] = 22'h 000000;  // +0.0000000000000000 = 2^ 2 * ln( 1 +  0 * 2^(- 2+1) + ( 0^2+ 0^2) * 2^(-2* 2) )   n =  2   d_n = 0 
assign u[4'b0000] [03] = 22'h 000000;  // +0.0000000000000000 = 2^ 3 * ln( 1 +  0 * 2^(- 3+1) + ( 0^2+ 0^2) * 2^(-2* 3) )   n =  3   d_n = 0 
assign u[4'b0000] [04] = 22'h 000000;  // +0.0000000000000000 = 2^ 4 * ln( 1 +  0 * 2^(- 4+1) + ( 0^2+ 0^2) * 2^(-2* 4) )   n =  4   d_n = 0 
assign u[4'b0000] [05] = 22'h 000000;  // +0.0000000000000000 = 2^ 5 * ln( 1 +  0 * 2^(- 5+1) + ( 0^2+ 0^2) * 2^(-2* 5) )   n =  5   d_n = 0 
assign u[4'b0000] [06] = 22'h 000000;  // +0.0000000000000000 = 2^ 6 * ln( 1 +  0 * 2^(- 6+1) + ( 0^2+ 0^2) * 2^(-2* 6) )   n =  6   d_n = 0 
assign u[4'b0000] [07] = 22'h 000000;  // +0.0000000000000000 = 2^ 7 * ln( 1 +  0 * 2^(- 7+1) + ( 0^2+ 0^2) * 2^(-2* 7) )   n =  7   d_n = 0 
assign u[4'b0000] [08] = 22'h 000000;  // +0.0000000000000000 = 2^ 8 * ln( 1 +  0 * 2^(- 8+1) + ( 0^2+ 0^2) * 2^(-2* 8) )   n =  8   d_n = 0 
assign u[4'b0000] [09] = 22'h 000000;  // +0.0000000000000000 = 2^ 9 * ln( 1 +  0 * 2^(- 9+1) + ( 0^2+ 0^2) * 2^(-2* 9) )   n =  9   d_n = 0 
assign u[4'b0000] [10] = 22'h 000000;  // +0.0000000000000000 = 2^10 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = 0 
assign u[4'b0000] [11] = 22'h 000000;  // +0.0000000000000000 = 2^11 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = 0 
assign u[4'b0000] [12] = 22'h 000000;  // +0.0000000000000000 = 2^12 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = 0 
assign u[4'b0000] [13] = 22'h 000000;  // +0.0000000000000000 = 2^13 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = 0 
assign u[4'b0000] [14] = 22'h 000000;  // +0.0000000000000000 = 2^14 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = 0 
assign u[4'b0000] [15] = 22'h 000000;  // +0.0000000000000000 = 2^15 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = 0 
assign u[4'b0000] [16] = 22'h 000000;  // +0.0000000000000000 = 2^16 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = 0 
assign u[4'b0000] [17] = 22'h 000000;  // +0.0000000000000000 = 2^17 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = 0 
assign u[4'b0000] [18] = 22'h 000000;  // +0.0000000000000000 = 2^18 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = 0 
assign u[4'b0000] [19] = 22'h 000000;  // +0.0000000000000000 = 2^19 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = 0 
assign u[4'b0000] [20] = 22'h 000000;  // +0.0000000000000000 = 2^20 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = 0 
assign u[4'b0000] [21] = 22'h 000000;  // +0.0000000000000000 = 2^21 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = 0 
assign u[4'b0000] [22] = 22'h 000000;  // +0.0000000000000000 = 2^22 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = 0 
assign u[4'b0000] [23] = 22'h 000000;  // +0.0000000000000000 = 2^23 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = 0 
assign u[4'b0000] [24] = 22'h 000000;  // +0.0000000000000000 = 2^24 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = 0 
assign u[4'b0000] [25] = 22'h 000000;  // +0.0000000000000000 = 2^25 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = 0 
assign u[4'b0000] [26] = 22'h 000000;  // +0.0000000000000000 = 2^26 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = 0 
assign u[4'b0000] [27] = 22'h 000000;  // +0.0000000000000000 = 2^27 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = 0 
assign u[4'b0000] [28] = 22'h 000000;  // +0.0000000000000000 = 2^28 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = 0 
assign u[4'b0000] [29] = 22'h 000000;  // +0.0000000000000000 = 2^29 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = 0 
assign u[4'b0000] [30] = 22'h 000000;  // +0.0000000000000000 = 2^30 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = 0 
assign u[4'b0000] [31] = 22'h 000000;  // +0.0000000000000000 = 2^31 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = 0 
assign u[4'b0000] [32] = 22'h 000000;  // +0.0000000000000000 = 2^32 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = 0 
assign u[4'b0000] [33] = 22'h 000000;  // +0.0000000000000000 = 2^33 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = 0 
assign u[4'b0000] [34] = 22'h 000000;  // +0.0000000000000000 = 2^34 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = 0 
assign u[4'b0000] [35] = 22'h 000000;  // +0.0000000000000000 = 2^35 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = 0 
assign u[4'b0000] [36] = 22'h 000000;  // +0.0000000000000000 = 2^36 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = 0 
assign u[4'b0000] [37] = 22'h 000000;  // +0.0000000000000000 = 2^37 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = 0 
assign u[4'b0000] [38] = 22'h 000000;  // +0.0000000000000000 = 2^38 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = 0 
assign u[4'b0000] [39] = 22'h 000000;  // +0.0000000000000000 = 2^39 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = 0 
assign u[4'b0000] [40] = 22'h 000000;  // +0.0000000000000000 = 2^40 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = 0 
assign u[4'b0000] [41] = 22'h 000000;  // +0.0000000000000000 = 2^41 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = 0 
assign u[4'b0000] [42] = 22'h 000000;  // +0.0000000000000000 = 2^42 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = 0 
assign u[4'b0000] [43] = 22'h 000000;  // +0.0000000000000000 = 2^43 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = 0 
assign u[4'b0000] [44] = 22'h 000000;  // +0.0000000000000000 = 2^44 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = 0 
assign u[4'b0000] [45] = 22'h 000000;  // +0.0000000000000000 = 2^45 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = 0 
assign u[4'b0000] [46] = 22'h 000000;  // +0.0000000000000000 = 2^46 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = 0 
assign u[4'b0000] [47] = 22'h 000000;  // +0.0000000000000000 = 2^47 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = 0 
assign u[4'b0000] [48] = 22'h 000000;  // +0.0000000000000000 = 2^48 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = 0 
assign u[4'b0000] [49] = 22'h 000000;  // +0.0000000000000000 = 2^49 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = 0 
assign u[4'b0000] [50] = 22'h 000000;  // +0.0000000000000000 = 2^50 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = 0 
assign u[4'b0000] [51] = 22'h 000000;  // +0.0000000000000000 = 2^51 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = 0 
assign u[4'b0000] [52] = 22'h 000000;  // +0.0000000000000000 = 2^52 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = 0 
assign u[4'b0000] [53] = 22'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = 0 
assign u[4'b0000] [54] = 22'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = 0 
assign u[4'b0000] [55] = 22'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = 0 
assign u[4'b0000] [56] = 22'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = 0 
assign u[4'b0000] [57] = 22'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = 0 
assign u[4'b0000] [58] = 22'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = 0 
assign u[4'b0000] [59] = 22'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = 0 
assign u[4'b0000] [60] = 22'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = 0 
assign u[4'b0000] [61] = 22'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = 0 
assign u[4'b0000] [62] = 22'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = 0 
assign u[4'b0000] [63] = 22'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = 0 
assign u[4'b0000] [64] = 22'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = 0 
assign u[4'b0001] [01] = 22'h 00019F;  // +1.6218604324326575 = 2^ 1 * ln( 1 +  1 * 2^(- 1+1) + ( 1^2+ 0^2) * 2^(-2* 1) )   n =  1   d_n = 1 
assign u[4'b0001] [02] = 22'h 0001C8;  // +1.7851484105136781 = 2^ 2 * ln( 1 +  1 * 2^(- 2+1) + ( 1^2+ 0^2) * 2^(-2* 2) )   n =  2   d_n = 1 
assign u[4'b0001] [03] = 22'h 0001E2;  // +1.8845285705021353 = 2^ 3 * ln( 1 +  1 * 2^(- 3+1) + ( 1^2+ 0^2) * 2^(-2* 3) )   n =  3   d_n = 1 
assign u[4'b0001] [04] = 22'h 0001F0;  // +1.9399878981259149 = 2^ 4 * ln( 1 +  1 * 2^(- 4+1) + ( 1^2+ 0^2) * 2^(-2* 4) )   n =  4   d_n = 1 
assign u[4'b0001] [05] = 22'h 0001F8;  // +1.9693861546722360 = 2^ 5 * ln( 1 +  1 * 2^(- 5+1) + ( 1^2+ 0^2) * 2^(-2* 5) )   n =  5   d_n = 1 
assign u[4'b0001] [06] = 22'h 0001FC;  // +1.9845358766035526 = 2^ 6 * ln( 1 +  1 * 2^(- 6+1) + ( 1^2+ 0^2) * 2^(-2* 6) )   n =  6   d_n = 1 
assign u[4'b0001] [07] = 22'h 0001FE;  // +1.9922279531660669 = 2^ 7 * ln( 1 +  1 * 2^(- 7+1) + ( 1^2+ 0^2) * 2^(-2* 7) )   n =  7   d_n = 1 
assign u[4'b0001] [08] = 22'h 0001FF;  // +1.9961038928165493 = 2^ 8 * ln( 1 +  1 * 2^(- 8+1) + ( 1^2+ 0^2) * 2^(-2* 8) )   n =  8   d_n = 1 
assign u[4'b0001] [09] = 22'h 0001FF;  // +1.9980494144120313 = 2^ 9 * ln( 1 +  1 * 2^(- 9+1) + ( 1^2+ 0^2) * 2^(-2* 9) )   n =  9   d_n = 1 
assign u[4'b0001] [10] = 22'h 0001FF;  // +1.9990240728175799 = 2^10 * ln( 1 +  1 * 2^(-10+1) + ( 1^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = 1 
assign u[4'b0001] [11] = 22'h 0001FF;  // +1.9995118776375345 = 2^11 * ln( 1 +  1 * 2^(-11+1) + ( 1^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = 1 
assign u[4'b0001] [12] = 22'h 0001FF;  // +1.9997558991041553 = 2^12 * ln( 1 +  1 * 2^(-12+1) + ( 1^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = 1 
assign u[4'b0001] [13] = 22'h 0001FF;  // +1.9998779396206980 = 2^13 * ln( 1 +  1 * 2^(-13+1) + ( 1^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = 1 
assign u[4'b0001] [14] = 22'h 0001FF;  // +1.9999389673271633 = 2^14 * ln( 1 +  1 * 2^(-14+1) + ( 1^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = 1 
assign u[4'b0001] [15] = 22'h 0001FF;  // +1.9999694830427426 = 2^15 * ln( 1 +  1 * 2^(-15+1) + ( 1^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = 1 
assign u[4'b0001] [16] = 22'h 0001FF;  // +1.9999847413661562 = 2^16 * ln( 1 +  1 * 2^(-16+1) + ( 1^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = 1 
assign u[4'b0001] [17] = 22'h 0001FF;  // +1.9999923706442737 = 2^17 * ln( 1 +  1 * 2^(-17+1) + ( 1^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = 1 
assign u[4'b0001] [18] = 22'h 0001FF;  // +1.9999961853124357 = 2^18 * ln( 1 +  1 * 2^(-18+1) + ( 1^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = 1 
assign u[4'b0001] [19] = 22'h 0001FF;  // +1.9999980926537926 = 2^19 * ln( 1 +  1 * 2^(-19+1) + ( 1^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = 1 
assign u[4'b0001] [20] = 22'h 0001FF;  // +1.9999990463262900 = 2^20 * ln( 1 +  1 * 2^(-20+1) + ( 1^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = 1 
assign u[4'b0001] [21] = 22'h 0001FF;  // +1.9999995231629935 = 2^21 * ln( 1 +  1 * 2^(-21+1) + ( 1^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = 1 
assign u[4'b0001] [22] = 22'h 0001FF;  // +1.9999997615814589 = 2^22 * ln( 1 +  1 * 2^(-22+1) + ( 1^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = 1 
assign u[4'b0001] [23] = 22'h 0001FF;  // +1.9999998807907200 = 2^23 * ln( 1 +  1 * 2^(-23+1) + ( 1^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = 1 
assign u[4'b0001] [24] = 22'h 0001FF;  // +1.9999999403953577 = 2^24 * ln( 1 +  1 * 2^(-24+1) + ( 1^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = 1 
assign u[4'b0001] [25] = 22'h 0001FF;  // +1.9999999701976783 = 2^25 * ln( 1 +  1 * 2^(-25+1) + ( 1^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = 1 
assign u[4'b0001] [26] = 22'h 0001FF;  // +1.9999999850988390 = 2^26 * ln( 1 +  1 * 2^(-26+1) + ( 1^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = 1 
assign u[4'b0001] [27] = 22'h 0001FF;  // +1.9999999925494194 = 2^27 * ln( 1 +  1 * 2^(-27+1) + ( 1^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = 1 
assign u[4'b0001] [28] = 22'h 0001FF;  // +1.9999999962747097 = 2^28 * ln( 1 +  1 * 2^(-28+1) + ( 1^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = 1 
assign u[4'b0001] [29] = 22'h 0001FF;  // +1.9999999981373549 = 2^29 * ln( 1 +  1 * 2^(-29+1) + ( 1^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = 1 
assign u[4'b0001] [30] = 22'h 0001FF;  // +1.9999999990686774 = 2^30 * ln( 1 +  1 * 2^(-30+1) + ( 1^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = 1 
assign u[4'b0001] [31] = 22'h 0001FF;  // +1.9999999995343387 = 2^31 * ln( 1 +  1 * 2^(-31+1) + ( 1^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = 1 
assign u[4'b0001] [32] = 22'h 0001FF;  // +1.9999999997671694 = 2^32 * ln( 1 +  1 * 2^(-32+1) + ( 1^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = 1 
assign u[4'b0001] [33] = 22'h 0001FF;  // +1.9999999998835847 = 2^33 * ln( 1 +  1 * 2^(-33+1) + ( 1^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = 1 
assign u[4'b0001] [34] = 22'h 0001FF;  // +1.9999999999417923 = 2^34 * ln( 1 +  1 * 2^(-34+1) + ( 1^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = 1 
assign u[4'b0001] [35] = 22'h 0001FF;  // +1.9999999999708962 = 2^35 * ln( 1 +  1 * 2^(-35+1) + ( 1^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = 1 
assign u[4'b0001] [36] = 22'h 0001FF;  // +1.9999999999854481 = 2^36 * ln( 1 +  1 * 2^(-36+1) + ( 1^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = 1 
assign u[4'b0001] [37] = 22'h 0001FF;  // +1.9999999999927240 = 2^37 * ln( 1 +  1 * 2^(-37+1) + ( 1^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = 1 
assign u[4'b0001] [38] = 22'h 0001FF;  // +1.9999999999963620 = 2^38 * ln( 1 +  1 * 2^(-38+1) + ( 1^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = 1 
assign u[4'b0001] [39] = 22'h 0001FF;  // +1.9999999999981810 = 2^39 * ln( 1 +  1 * 2^(-39+1) + ( 1^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = 1 
assign u[4'b0001] [40] = 22'h 0001FF;  // +1.9999999999990905 = 2^40 * ln( 1 +  1 * 2^(-40+1) + ( 1^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = 1 
assign u[4'b0001] [41] = 22'h 0001FF;  // +1.9999999999995453 = 2^41 * ln( 1 +  1 * 2^(-41+1) + ( 1^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = 1 
assign u[4'b0001] [42] = 22'h 0001FF;  // +1.9999999999997726 = 2^42 * ln( 1 +  1 * 2^(-42+1) + ( 1^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = 1 
assign u[4'b0001] [43] = 22'h 0001FF;  // +1.9999999999998863 = 2^43 * ln( 1 +  1 * 2^(-43+1) + ( 1^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = 1 
assign u[4'b0001] [44] = 22'h 0001FF;  // +1.9999999999999432 = 2^44 * ln( 1 +  1 * 2^(-44+1) + ( 1^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = 1 
assign u[4'b0001] [45] = 22'h 0001FF;  // +1.9999999999999716 = 2^45 * ln( 1 +  1 * 2^(-45+1) + ( 1^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = 1 
assign u[4'b0001] [46] = 22'h 0001FF;  // +1.9999999999999858 = 2^46 * ln( 1 +  1 * 2^(-46+1) + ( 1^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = 1 
assign u[4'b0001] [47] = 22'h 0001FF;  // +1.9999999999999929 = 2^47 * ln( 1 +  1 * 2^(-47+1) + ( 1^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = 1 
assign u[4'b0001] [48] = 22'h 0001FF;  // +1.9999999999999964 = 2^48 * ln( 1 +  1 * 2^(-48+1) + ( 1^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = 1 
assign u[4'b0001] [49] = 22'h 0001FF;  // +1.9999999999999982 = 2^49 * ln( 1 +  1 * 2^(-49+1) + ( 1^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = 1 
assign u[4'b0001] [50] = 22'h 0001FF;  // +1.9999999999999991 = 2^50 * ln( 1 +  1 * 2^(-50+1) + ( 1^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = 1 
assign u[4'b0001] [51] = 22'h 0001FF;  // +1.9999999999999996 = 2^51 * ln( 1 +  1 * 2^(-51+1) + ( 1^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = 1 
assign u[4'b0001] [52] = 22'h 0001FF;  // +1.9999999999999998 = 2^52 * ln( 1 +  1 * 2^(-52+1) + ( 1^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = 1 
assign u[4'b0001] [53] = 22'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  1 * 2^(-53+1) + ( 1^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = 1 
assign u[4'b0001] [54] = 22'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  1 * 2^(-54+1) + ( 1^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = 1 
assign u[4'b0001] [55] = 22'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  1 * 2^(-55+1) + ( 1^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = 1 
assign u[4'b0001] [56] = 22'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  1 * 2^(-56+1) + ( 1^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = 1 
assign u[4'b0001] [57] = 22'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  1 * 2^(-57+1) + ( 1^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = 1 
assign u[4'b0001] [58] = 22'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  1 * 2^(-58+1) + ( 1^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = 1 
assign u[4'b0001] [59] = 22'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  1 * 2^(-59+1) + ( 1^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = 1 
assign u[4'b0001] [60] = 22'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  1 * 2^(-60+1) + ( 1^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = 1 
assign u[4'b0001] [61] = 22'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  1 * 2^(-61+1) + ( 1^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = 1 
assign u[4'b0001] [62] = 22'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  1 * 2^(-62+1) + ( 1^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = 1 
assign u[4'b0001] [63] = 22'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  1 * 2^(-63+1) + ( 1^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = 1 
assign u[4'b0001] [64] = 22'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  1 * 2^(-64+1) + ( 1^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = 1 
assign u[4'b0010] [01] = 22'h 000000;  // +0.0000000000000000 = 2^ 1 * ln( 1 +  0 * 2^(- 1+1) + ( 0^2+ 0^2) * 2^(-2* 1) )   n =  1   d_n = -0 
assign u[4'b0010] [02] = 22'h 000000;  // +0.0000000000000000 = 2^ 2 * ln( 1 +  0 * 2^(- 2+1) + ( 0^2+ 0^2) * 2^(-2* 2) )   n =  2   d_n = -0 
assign u[4'b0010] [03] = 22'h 000000;  // +0.0000000000000000 = 2^ 3 * ln( 1 +  0 * 2^(- 3+1) + ( 0^2+ 0^2) * 2^(-2* 3) )   n =  3   d_n = -0 
assign u[4'b0010] [04] = 22'h 000000;  // +0.0000000000000000 = 2^ 4 * ln( 1 +  0 * 2^(- 4+1) + ( 0^2+ 0^2) * 2^(-2* 4) )   n =  4   d_n = -0 
assign u[4'b0010] [05] = 22'h 000000;  // +0.0000000000000000 = 2^ 5 * ln( 1 +  0 * 2^(- 5+1) + ( 0^2+ 0^2) * 2^(-2* 5) )   n =  5   d_n = -0 
assign u[4'b0010] [06] = 22'h 000000;  // +0.0000000000000000 = 2^ 6 * ln( 1 +  0 * 2^(- 6+1) + ( 0^2+ 0^2) * 2^(-2* 6) )   n =  6   d_n = -0 
assign u[4'b0010] [07] = 22'h 000000;  // +0.0000000000000000 = 2^ 7 * ln( 1 +  0 * 2^(- 7+1) + ( 0^2+ 0^2) * 2^(-2* 7) )   n =  7   d_n = -0 
assign u[4'b0010] [08] = 22'h 000000;  // +0.0000000000000000 = 2^ 8 * ln( 1 +  0 * 2^(- 8+1) + ( 0^2+ 0^2) * 2^(-2* 8) )   n =  8   d_n = -0 
assign u[4'b0010] [09] = 22'h 000000;  // +0.0000000000000000 = 2^ 9 * ln( 1 +  0 * 2^(- 9+1) + ( 0^2+ 0^2) * 2^(-2* 9) )   n =  9   d_n = -0 
assign u[4'b0010] [10] = 22'h 000000;  // +0.0000000000000000 = 2^10 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = -0 
assign u[4'b0010] [11] = 22'h 000000;  // +0.0000000000000000 = 2^11 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = -0 
assign u[4'b0010] [12] = 22'h 000000;  // +0.0000000000000000 = 2^12 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = -0 
assign u[4'b0010] [13] = 22'h 000000;  // +0.0000000000000000 = 2^13 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = -0 
assign u[4'b0010] [14] = 22'h 000000;  // +0.0000000000000000 = 2^14 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = -0 
assign u[4'b0010] [15] = 22'h 000000;  // +0.0000000000000000 = 2^15 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = -0 
assign u[4'b0010] [16] = 22'h 000000;  // +0.0000000000000000 = 2^16 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = -0 
assign u[4'b0010] [17] = 22'h 000000;  // +0.0000000000000000 = 2^17 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = -0 
assign u[4'b0010] [18] = 22'h 000000;  // +0.0000000000000000 = 2^18 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = -0 
assign u[4'b0010] [19] = 22'h 000000;  // +0.0000000000000000 = 2^19 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = -0 
assign u[4'b0010] [20] = 22'h 000000;  // +0.0000000000000000 = 2^20 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = -0 
assign u[4'b0010] [21] = 22'h 000000;  // +0.0000000000000000 = 2^21 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = -0 
assign u[4'b0010] [22] = 22'h 000000;  // +0.0000000000000000 = 2^22 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = -0 
assign u[4'b0010] [23] = 22'h 000000;  // +0.0000000000000000 = 2^23 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = -0 
assign u[4'b0010] [24] = 22'h 000000;  // +0.0000000000000000 = 2^24 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = -0 
assign u[4'b0010] [25] = 22'h 000000;  // +0.0000000000000000 = 2^25 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = -0 
assign u[4'b0010] [26] = 22'h 000000;  // +0.0000000000000000 = 2^26 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = -0 
assign u[4'b0010] [27] = 22'h 000000;  // +0.0000000000000000 = 2^27 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = -0 
assign u[4'b0010] [28] = 22'h 000000;  // +0.0000000000000000 = 2^28 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = -0 
assign u[4'b0010] [29] = 22'h 000000;  // +0.0000000000000000 = 2^29 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = -0 
assign u[4'b0010] [30] = 22'h 000000;  // +0.0000000000000000 = 2^30 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = -0 
assign u[4'b0010] [31] = 22'h 000000;  // +0.0000000000000000 = 2^31 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = -0 
assign u[4'b0010] [32] = 22'h 000000;  // +0.0000000000000000 = 2^32 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = -0 
assign u[4'b0010] [33] = 22'h 000000;  // +0.0000000000000000 = 2^33 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = -0 
assign u[4'b0010] [34] = 22'h 000000;  // +0.0000000000000000 = 2^34 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = -0 
assign u[4'b0010] [35] = 22'h 000000;  // +0.0000000000000000 = 2^35 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = -0 
assign u[4'b0010] [36] = 22'h 000000;  // +0.0000000000000000 = 2^36 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = -0 
assign u[4'b0010] [37] = 22'h 000000;  // +0.0000000000000000 = 2^37 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = -0 
assign u[4'b0010] [38] = 22'h 000000;  // +0.0000000000000000 = 2^38 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = -0 
assign u[4'b0010] [39] = 22'h 000000;  // +0.0000000000000000 = 2^39 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = -0 
assign u[4'b0010] [40] = 22'h 000000;  // +0.0000000000000000 = 2^40 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = -0 
assign u[4'b0010] [41] = 22'h 000000;  // +0.0000000000000000 = 2^41 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = -0 
assign u[4'b0010] [42] = 22'h 000000;  // +0.0000000000000000 = 2^42 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = -0 
assign u[4'b0010] [43] = 22'h 000000;  // +0.0000000000000000 = 2^43 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = -0 
assign u[4'b0010] [44] = 22'h 000000;  // +0.0000000000000000 = 2^44 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = -0 
assign u[4'b0010] [45] = 22'h 000000;  // +0.0000000000000000 = 2^45 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = -0 
assign u[4'b0010] [46] = 22'h 000000;  // +0.0000000000000000 = 2^46 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = -0 
assign u[4'b0010] [47] = 22'h 000000;  // +0.0000000000000000 = 2^47 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = -0 
assign u[4'b0010] [48] = 22'h 000000;  // +0.0000000000000000 = 2^48 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = -0 
assign u[4'b0010] [49] = 22'h 000000;  // +0.0000000000000000 = 2^49 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = -0 
assign u[4'b0010] [50] = 22'h 000000;  // +0.0000000000000000 = 2^50 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = -0 
assign u[4'b0010] [51] = 22'h 000000;  // +0.0000000000000000 = 2^51 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = -0 
assign u[4'b0010] [52] = 22'h 000000;  // +0.0000000000000000 = 2^52 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = -0 
assign u[4'b0010] [53] = 22'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = -0 
assign u[4'b0010] [54] = 22'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = -0 
assign u[4'b0010] [55] = 22'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = -0 
assign u[4'b0010] [56] = 22'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = -0 
assign u[4'b0010] [57] = 22'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = -0 
assign u[4'b0010] [58] = 22'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = -0 
assign u[4'b0010] [59] = 22'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = -0 
assign u[4'b0010] [60] = 22'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = -0 
assign u[4'b0010] [61] = 22'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = -0 
assign u[4'b0010] [62] = 22'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = -0 
assign u[4'b0010] [63] = 22'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = -0 
assign u[4'b0010] [64] = 22'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = -0 
assign u[4'b0011] [01] = 22'h 3FFD3A;  // -2.7725887222397811 = 2^ 1 * ln( 1 + -1 * 2^(- 1+1) + (-1^2+ 0^2) * 2^(-2* 1) )   n =  1   d_n = -1 
assign u[4'b0011] [02] = 22'h 3FFDB2;  // -2.3014565796142472 = 2^ 2 * ln( 1 + -1 * 2^(- 2+1) + (-1^2+ 0^2) * 2^(-2* 2) )   n =  2   d_n = -1 
assign u[4'b0011] [03] = 22'h 3FFDDD;  // -2.1365022819923620 = 2^ 3 * ln( 1 + -1 * 2^(- 3+1) + (-1^2+ 0^2) * 2^(-2* 3) )   n =  3   d_n = -1 
assign u[4'b0011] [04] = 22'h 3FFDEF;  // -2.0652326764022777 = 2^ 4 * ln( 1 + -1 * 2^(- 4+1) + (-1^2+ 0^2) * 2^(-2* 4) )   n =  4   d_n = -1 
assign u[4'b0011] [05] = 22'h 3FFDF7;  // -2.0319166921331391 = 2^ 5 * ln( 1 + -1 * 2^(- 5+1) + (-1^2+ 0^2) * 2^(-2* 5) )   n =  5   d_n = -1 
assign u[4'b0011] [06] = 22'h 3FFDFB;  // -2.0157896919218135 = 2^ 6 * ln( 1 + -1 * 2^(- 6+1) + (-1^2+ 0^2) * 2^(-2* 6) )   n =  6   d_n = -1 
assign u[4'b0011] [07] = 22'h 3FFDFD;  // -2.0078534300226285 = 2^ 7 * ln( 1 + -1 * 2^(- 7+1) + (-1^2+ 0^2) * 2^(-2* 7) )   n =  7   d_n = -1 
assign u[4'b0011] [08] = 22'h 3FFDFE;  // -2.0039164524218003 = 2^ 8 * ln( 1 + -1 * 2^(- 8+1) + (-1^2+ 0^2) * 2^(-2* 8) )   n =  8   d_n = -1 
assign u[4'b0011] [09] = 22'h 3FFDFF;  // -2.0019556718626310 = 2^ 9 * ln( 1 + -1 * 2^(- 9+1) + (-1^2+ 0^2) * 2^(-2* 9) )   n =  9   d_n = -1 
assign u[4'b0011] [10] = 22'h 3FFDFF;  // -2.0009771987489029 = 2^10 * ln( 1 + -1 * 2^(-10+1) + (-1^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = -1 
assign u[4'b0011] [11] = 22'h 3FFDFF;  // -2.0004884402539500 = 2^11 * ln( 1 + -1 * 2^(-11+1) + (-1^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = -1 
assign u[4'b0011] [12] = 22'h 3FFDFF;  // -2.0002441803687074 = 2^12 * ln( 1 + -1 * 2^(-12+1) + (-1^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = -1 
assign u[4'b0011] [13] = 22'h 3FFDFF;  // -2.0001220802475173 = 2^13 * ln( 1 + -1 * 2^(-13+1) + (-1^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = -1 
assign u[4'b0011] [14] = 22'h 3FFDFF;  // -2.0000610376398904 = 2^14 * ln( 1 + -1 * 2^(-14+1) + (-1^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = -1 
assign u[4'b0011] [15] = 22'h 3FFDFF;  // -2.0000305181990208 = 2^15 * ln( 1 + -1 * 2^(-15+1) + (-1^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = -1 
assign u[4'b0011] [16] = 22'h 3FFDFF;  // -2.0000152589442846 = 2^16 * ln( 1 + -1 * 2^(-16+1) + (-1^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = -1 
assign u[4'b0011] [17] = 22'h 3FFDFF;  // -2.0000076294333367 = 2^17 * ln( 1 + -1 * 2^(-17+1) + (-1^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = -1 
assign u[4'b0011] [18] = 22'h 3FFDFF;  // -2.0000038147069668 = 2^18 * ln( 1 + -1 * 2^(-18+1) + (-1^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = -1 
assign u[4'b0011] [19] = 22'h 3FFDFF;  // -2.0000019073510580 = 2^19 * ln( 1 + -1 * 2^(-19+1) + (-1^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = -1 
assign u[4'b0011] [20] = 22'h 3FFDFF;  // -2.0000009536749226 = 2^20 * ln( 1 + -1 * 2^(-20+1) + (-1^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = -1 
assign u[4'b0011] [21] = 22'h 3FFDFF;  // -2.0000004768373096 = 2^21 * ln( 1 + -1 * 2^(-21+1) + (-1^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = -1 
assign u[4'b0011] [22] = 22'h 3FFDFF;  // -2.0000002384186168 = 2^22 * ln( 1 + -1 * 2^(-22+1) + (-1^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = -1 
assign u[4'b0011] [23] = 22'h 3FFDFF;  // -2.0000001192092989 = 2^23 * ln( 1 + -1 * 2^(-23+1) + (-1^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = -1 
assign u[4'b0011] [24] = 22'h 3FFDFF;  // -2.0000000596046470 = 2^24 * ln( 1 + -1 * 2^(-24+1) + (-1^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = -1 
assign u[4'b0011] [25] = 22'h 3FFDFF;  // -2.0000000298023228 = 2^25 * ln( 1 + -1 * 2^(-25+1) + (-1^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = -1 
assign u[4'b0011] [26] = 22'h 3FFDFF;  // -2.0000000149011612 = 2^26 * ln( 1 + -1 * 2^(-26+1) + (-1^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = -1 
assign u[4'b0011] [27] = 22'h 3FFDFF;  // -2.0000000074505806 = 2^27 * ln( 1 + -1 * 2^(-27+1) + (-1^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = -1 
assign u[4'b0011] [28] = 22'h 3FFDFF;  // -2.0000000037252903 = 2^28 * ln( 1 + -1 * 2^(-28+1) + (-1^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = -1 
assign u[4'b0011] [29] = 22'h 3FFDFF;  // -2.0000000018626451 = 2^29 * ln( 1 + -1 * 2^(-29+1) + (-1^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = -1 
assign u[4'b0011] [30] = 22'h 3FFDFF;  // -2.0000000009313226 = 2^30 * ln( 1 + -1 * 2^(-30+1) + (-1^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = -1 
assign u[4'b0011] [31] = 22'h 3FFDFF;  // -2.0000000004656613 = 2^31 * ln( 1 + -1 * 2^(-31+1) + (-1^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = -1 
assign u[4'b0011] [32] = 22'h 3FFDFF;  // -2.0000000002328306 = 2^32 * ln( 1 + -1 * 2^(-32+1) + (-1^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = -1 
assign u[4'b0011] [33] = 22'h 3FFDFF;  // -2.0000000001164153 = 2^33 * ln( 1 + -1 * 2^(-33+1) + (-1^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = -1 
assign u[4'b0011] [34] = 22'h 3FFDFF;  // -2.0000000000582077 = 2^34 * ln( 1 + -1 * 2^(-34+1) + (-1^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = -1 
assign u[4'b0011] [35] = 22'h 3FFDFF;  // -2.0000000000291038 = 2^35 * ln( 1 + -1 * 2^(-35+1) + (-1^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = -1 
assign u[4'b0011] [36] = 22'h 3FFDFF;  // -2.0000000000145519 = 2^36 * ln( 1 + -1 * 2^(-36+1) + (-1^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = -1 
assign u[4'b0011] [37] = 22'h 3FFDFF;  // -2.0000000000072760 = 2^37 * ln( 1 + -1 * 2^(-37+1) + (-1^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = -1 
assign u[4'b0011] [38] = 22'h 3FFDFF;  // -2.0000000000036380 = 2^38 * ln( 1 + -1 * 2^(-38+1) + (-1^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = -1 
assign u[4'b0011] [39] = 22'h 3FFDFF;  // -2.0000000000018190 = 2^39 * ln( 1 + -1 * 2^(-39+1) + (-1^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = -1 
assign u[4'b0011] [40] = 22'h 3FFE00;  // -2.0000000000009095 = 2^40 * ln( 1 + -1 * 2^(-40+1) + (-1^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = -1 
assign u[4'b0011] [41] = 22'h 3FFE00;  // -2.0000000000004547 = 2^41 * ln( 1 + -1 * 2^(-41+1) + (-1^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = -1 
assign u[4'b0011] [42] = 22'h 3FFE00;  // -2.0000000000002274 = 2^42 * ln( 1 + -1 * 2^(-42+1) + (-1^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = -1 
assign u[4'b0011] [43] = 22'h 3FFE00;  // -2.0000000000001137 = 2^43 * ln( 1 + -1 * 2^(-43+1) + (-1^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = -1 
assign u[4'b0011] [44] = 22'h 3FFE00;  // -2.0000000000000568 = 2^44 * ln( 1 + -1 * 2^(-44+1) + (-1^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = -1 
assign u[4'b0011] [45] = 22'h 3FFE00;  // -2.0000000000000284 = 2^45 * ln( 1 + -1 * 2^(-45+1) + (-1^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = -1 
assign u[4'b0011] [46] = 22'h 3FFE00;  // -2.0000000000000142 = 2^46 * ln( 1 + -1 * 2^(-46+1) + (-1^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = -1 
assign u[4'b0011] [47] = 22'h 3FFE00;  // -2.0000000000000071 = 2^47 * ln( 1 + -1 * 2^(-47+1) + (-1^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = -1 
assign u[4'b0011] [48] = 22'h 3FFE00;  // -2.0000000000000036 = 2^48 * ln( 1 + -1 * 2^(-48+1) + (-1^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = -1 
assign u[4'b0011] [49] = 22'h 3FFE00;  // -2.0000000000000018 = 2^49 * ln( 1 + -1 * 2^(-49+1) + (-1^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = -1 
assign u[4'b0011] [50] = 22'h 3FFE00;  // -2.0000000000000009 = 2^50 * ln( 1 + -1 * 2^(-50+1) + (-1^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = -1 
assign u[4'b0011] [51] = 22'h 3FFE00;  // -2.0000000000000004 = 2^51 * ln( 1 + -1 * 2^(-51+1) + (-1^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = -1 
assign u[4'b0011] [52] = 22'h 3FFE00;  // -2.0000000000000004 = 2^52 * ln( 1 + -1 * 2^(-52+1) + (-1^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = -1 
assign u[4'b0011] [53] = 22'h 3FFE00;  // -2.0000000000000000 = 2^53 * ln( 1 + -1 * 2^(-53+1) + (-1^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = -1 
assign u[4'b0011] [54] = 22'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 + -1 * 2^(-54+1) + (-1^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = -1 
assign u[4'b0011] [55] = 22'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 + -1 * 2^(-55+1) + (-1^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = -1 
assign u[4'b0011] [56] = 22'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 + -1 * 2^(-56+1) + (-1^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = -1 
assign u[4'b0011] [57] = 22'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 + -1 * 2^(-57+1) + (-1^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = -1 
assign u[4'b0011] [58] = 22'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 + -1 * 2^(-58+1) + (-1^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = -1 
assign u[4'b0011] [59] = 22'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 + -1 * 2^(-59+1) + (-1^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = -1 
assign u[4'b0011] [60] = 22'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 + -1 * 2^(-60+1) + (-1^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = -1 
assign u[4'b0011] [61] = 22'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 + -1 * 2^(-61+1) + (-1^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = -1 
assign u[4'b0011] [62] = 22'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 + -1 * 2^(-62+1) + (-1^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = -1 
assign u[4'b0011] [63] = 22'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 + -1 * 2^(-63+1) + (-1^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = -1 
assign u[4'b0011] [64] = 22'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 + -1 * 2^(-64+1) + (-1^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = -1 
assign u[4'b0100] [01] = 22'h 000072;  // +0.4462871026284197 = 2^ 1 * ln( 1 +  0 * 2^(- 1+1) + ( 0^2+ 1^2) * 2^(-2* 1) )   n =  1   d_n = 0+1i 
assign u[4'b0100] [02] = 22'h 00003E;  // +0.2424984872657394 = 2^ 2 * ln( 1 +  0 * 2^(- 2+1) + ( 0^2+ 1^2) * 2^(-2* 2) )   n =  2   d_n = 0+1i 
assign u[4'b0100] [03] = 22'h 00001F;  // +0.1240334922877210 = 2^ 3 * ln( 1 +  0 * 2^(- 3+1) + ( 0^2+ 1^2) * 2^(-2* 3) )   n =  3   d_n = 0+1i 
assign u[4'b0100] [04] = 22'h 00000F;  // +0.0623782466505195 = 2^ 4 * ln( 1 +  0 * 2^(- 4+1) + ( 0^2+ 1^2) * 2^(-2* 4) )   n =  4   d_n = 0+1i 
assign u[4'b0100] [05] = 22'h 000007;  // +0.0312347511377731 = 2^ 5 * ln( 1 +  0 * 2^(- 5+1) + ( 0^2+ 1^2) * 2^(-2* 5) )   n =  5   d_n = 0+1i 
assign u[4'b0100] [06] = 22'h 000003;  // +0.0156230929617406 = 2^ 6 * ln( 1 +  0 * 2^(- 6+1) + ( 0^2+ 1^2) * 2^(-2* 6) )   n =  6   d_n = 0+1i 
assign u[4'b0100] [07] = 22'h 000001;  // +0.0078122615911219 = 2^ 7 * ln( 1 +  0 * 2^(- 7+1) + ( 0^2+ 1^2) * 2^(-2* 7) )   n =  7   d_n = 0+1i 
assign u[4'b0100] [08] = 22'h 000000;  // +0.0039062201979808 = 2^ 8 * ln( 1 +  0 * 2^(- 8+1) + ( 0^2+ 1^2) * 2^(-2* 8) )   n =  8   d_n = 0+1i 
assign u[4'b0100] [09] = 22'h 000000;  // +0.0019531212747156 = 2^ 9 * ln( 1 +  0 * 2^(- 9+1) + ( 0^2+ 1^2) * 2^(-2* 9) )   n =  9   d_n = 0+1i 
assign u[4'b0100] [10] = 22'h 000000;  // +0.0009765620343389 = 2^10 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 1^2) * 2^(-2*10) )   n = 10   d_n = 0+1i 
assign u[4'b0100] [11] = 22'h 000000;  // +0.0004882811917923 = 2^11 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 1^2) * 2^(-2*11) )   n = 11   d_n = 0+1i 
assign u[4'b0100] [12] = 22'h 000000;  // +0.0002441406177240 = 2^12 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 1^2) * 2^(-2*12) )   n = 12   d_n = 0+1i 
assign u[4'b0100] [13] = 22'h 000000;  // +0.0001220703120453 = 2^13 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 1^2) * 2^(-2*13) )   n = 13   d_n = 0+1i 
assign u[4'b0100] [14] = 22'h 000000;  // +0.0000610351561932 = 2^14 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 1^2) * 2^(-2*14) )   n = 14   d_n = 0+1i 
assign u[4'b0100] [15] = 22'h 000000;  // +0.0000305175781179 = 2^15 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 1^2) * 2^(-2*15) )   n = 15   d_n = 0+1i 
assign u[4'b0100] [16] = 22'h 000000;  // +0.0000152587890616 = 2^16 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 1^2) * 2^(-2*16) )   n = 16   d_n = 0+1i 
assign u[4'b0100] [17] = 22'h 000000;  // +0.0000076293945311 = 2^17 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 1^2) * 2^(-2*17) )   n = 17   d_n = 0+1i 
assign u[4'b0100] [18] = 22'h 000000;  // +0.0000038146972656 = 2^18 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 1^2) * 2^(-2*18) )   n = 18   d_n = 0+1i 
assign u[4'b0100] [19] = 22'h 000000;  // +0.0000019073486328 = 2^19 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 1^2) * 2^(-2*19) )   n = 19   d_n = 0+1i 
assign u[4'b0100] [20] = 22'h 000000;  // +0.0000009536743164 = 2^20 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 1^2) * 2^(-2*20) )   n = 20   d_n = 0+1i 
assign u[4'b0100] [21] = 22'h 000000;  // +0.0000004768371582 = 2^21 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 1^2) * 2^(-2*21) )   n = 21   d_n = 0+1i 
assign u[4'b0100] [22] = 22'h 000000;  // +0.0000002384185791 = 2^22 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 1^2) * 2^(-2*22) )   n = 22   d_n = 0+1i 
assign u[4'b0100] [23] = 22'h 000000;  // +0.0000001192092896 = 2^23 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 1^2) * 2^(-2*23) )   n = 23   d_n = 0+1i 
assign u[4'b0100] [24] = 22'h 000000;  // +0.0000000596046448 = 2^24 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 1^2) * 2^(-2*24) )   n = 24   d_n = 0+1i 
assign u[4'b0100] [25] = 22'h 000000;  // +0.0000000298023224 = 2^25 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 1^2) * 2^(-2*25) )   n = 25   d_n = 0+1i 
assign u[4'b0100] [26] = 22'h 000000;  // +0.0000000000000000 = 2^26 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 1^2) * 2^(-2*26) )   n = 26   d_n = 0+1i 
assign u[4'b0100] [27] = 22'h 000000;  // +0.0000000000000000 = 2^27 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 1^2) * 2^(-2*27) )   n = 27   d_n = 0+1i 
assign u[4'b0100] [28] = 22'h 000000;  // +0.0000000000000000 = 2^28 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 1^2) * 2^(-2*28) )   n = 28   d_n = 0+1i 
assign u[4'b0100] [29] = 22'h 000000;  // +0.0000000000000000 = 2^29 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 1^2) * 2^(-2*29) )   n = 29   d_n = 0+1i 
assign u[4'b0100] [30] = 22'h 000000;  // +0.0000000000000000 = 2^30 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 1^2) * 2^(-2*30) )   n = 30   d_n = 0+1i 
assign u[4'b0100] [31] = 22'h 000000;  // +0.0000000000000000 = 2^31 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 1^2) * 2^(-2*31) )   n = 31   d_n = 0+1i 
assign u[4'b0100] [32] = 22'h 000000;  // +0.0000000000000000 = 2^32 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 1^2) * 2^(-2*32) )   n = 32   d_n = 0+1i 
assign u[4'b0100] [33] = 22'h 000000;  // +0.0000000000000000 = 2^33 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 1^2) * 2^(-2*33) )   n = 33   d_n = 0+1i 
assign u[4'b0100] [34] = 22'h 000000;  // +0.0000000000000000 = 2^34 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 1^2) * 2^(-2*34) )   n = 34   d_n = 0+1i 
assign u[4'b0100] [35] = 22'h 000000;  // +0.0000000000000000 = 2^35 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 1^2) * 2^(-2*35) )   n = 35   d_n = 0+1i 
assign u[4'b0100] [36] = 22'h 000000;  // +0.0000000000000000 = 2^36 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 1^2) * 2^(-2*36) )   n = 36   d_n = 0+1i 
assign u[4'b0100] [37] = 22'h 000000;  // +0.0000000000000000 = 2^37 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 1^2) * 2^(-2*37) )   n = 37   d_n = 0+1i 
assign u[4'b0100] [38] = 22'h 000000;  // +0.0000000000000000 = 2^38 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 1^2) * 2^(-2*38) )   n = 38   d_n = 0+1i 
assign u[4'b0100] [39] = 22'h 000000;  // +0.0000000000000000 = 2^39 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 1^2) * 2^(-2*39) )   n = 39   d_n = 0+1i 
assign u[4'b0100] [40] = 22'h 000000;  // +0.0000000000000000 = 2^40 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 1^2) * 2^(-2*40) )   n = 40   d_n = 0+1i 
assign u[4'b0100] [41] = 22'h 000000;  // +0.0000000000000000 = 2^41 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 1^2) * 2^(-2*41) )   n = 41   d_n = 0+1i 
assign u[4'b0100] [42] = 22'h 000000;  // +0.0000000000000000 = 2^42 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 1^2) * 2^(-2*42) )   n = 42   d_n = 0+1i 
assign u[4'b0100] [43] = 22'h 000000;  // +0.0000000000000000 = 2^43 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 1^2) * 2^(-2*43) )   n = 43   d_n = 0+1i 
assign u[4'b0100] [44] = 22'h 000000;  // +0.0000000000000000 = 2^44 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 1^2) * 2^(-2*44) )   n = 44   d_n = 0+1i 
assign u[4'b0100] [45] = 22'h 000000;  // +0.0000000000000000 = 2^45 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 1^2) * 2^(-2*45) )   n = 45   d_n = 0+1i 
assign u[4'b0100] [46] = 22'h 000000;  // +0.0000000000000000 = 2^46 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 1^2) * 2^(-2*46) )   n = 46   d_n = 0+1i 
assign u[4'b0100] [47] = 22'h 000000;  // +0.0000000000000000 = 2^47 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 1^2) * 2^(-2*47) )   n = 47   d_n = 0+1i 
assign u[4'b0100] [48] = 22'h 000000;  // +0.0000000000000000 = 2^48 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 1^2) * 2^(-2*48) )   n = 48   d_n = 0+1i 
assign u[4'b0100] [49] = 22'h 000000;  // +0.0000000000000000 = 2^49 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 1^2) * 2^(-2*49) )   n = 49   d_n = 0+1i 
assign u[4'b0100] [50] = 22'h 000000;  // +0.0000000000000000 = 2^50 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 1^2) * 2^(-2*50) )   n = 50   d_n = 0+1i 
assign u[4'b0100] [51] = 22'h 000000;  // +0.0000000000000000 = 2^51 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 1^2) * 2^(-2*51) )   n = 51   d_n = 0+1i 
assign u[4'b0100] [52] = 22'h 000000;  // +0.0000000000000000 = 2^52 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 1^2) * 2^(-2*52) )   n = 52   d_n = 0+1i 
assign u[4'b0100] [53] = 22'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 1^2) * 2^(-2*53) )   n = 53   d_n = 0+1i 
assign u[4'b0100] [54] = 22'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 1^2) * 2^(-2*54) )   n = 54   d_n = 0+1i 
assign u[4'b0100] [55] = 22'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 1^2) * 2^(-2*55) )   n = 55   d_n = 0+1i 
assign u[4'b0100] [56] = 22'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 1^2) * 2^(-2*56) )   n = 56   d_n = 0+1i 
assign u[4'b0100] [57] = 22'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 1^2) * 2^(-2*57) )   n = 57   d_n = 0+1i 
assign u[4'b0100] [58] = 22'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 1^2) * 2^(-2*58) )   n = 58   d_n = 0+1i 
assign u[4'b0100] [59] = 22'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 1^2) * 2^(-2*59) )   n = 59   d_n = 0+1i 
assign u[4'b0100] [60] = 22'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 1^2) * 2^(-2*60) )   n = 60   d_n = 0+1i 
assign u[4'b0100] [61] = 22'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 1^2) * 2^(-2*61) )   n = 61   d_n = 0+1i 
assign u[4'b0100] [62] = 22'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 1^2) * 2^(-2*62) )   n = 62   d_n = 0+1i 
assign u[4'b0100] [63] = 22'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 1^2) * 2^(-2*63) )   n = 63   d_n = 0+1i 
assign u[4'b0100] [64] = 22'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 1^2) * 2^(-2*64) )   n = 64   d_n = 0+1i 
assign u[4'b0101] [01] = 22'h 0001D5;  // +1.8325814637483104 = 2^ 1 * ln( 1 +  1 * 2^(- 1+1) + ( 1^2+ 1^2) * 2^(-2* 1) )   n =  1   d_n = 1+1i 
assign u[4'b0101] [02] = 22'h 0001F1;  // +1.9420312631268026 = 2^ 2 * ln( 1 +  1 * 2^(- 2+1) + ( 1^2+ 1^2) * 2^(-2* 2) )   n =  2   d_n = 1+1i 
assign u[4'b0101] [03] = 22'h 0001FB;  // +1.9826893112366513 = 2^ 3 * ln( 1 +  1 * 2^(- 3+1) + ( 1^2+ 1^2) * 2^(-2* 3) )   n =  3   d_n = 1+1i 
assign u[4'b0101] [04] = 22'h 0001FE;  // +1.9952556560153185 = 2^ 4 * ln( 1 +  1 * 2^(- 4+1) + ( 1^2+ 1^2) * 2^(-2* 4) )   n =  4   d_n = 1+1i 
assign u[4'b0101] [05] = 22'h 0001FF;  // +1.9987574279595595 = 2^ 5 * ln( 1 +  1 * 2^(- 5+1) + ( 1^2+ 1^2) * 2^(-2* 5) )   n =  5   d_n = 1+1i 
assign u[4'b0101] [06] = 22'h 0001FF;  // +1.9996820132261188 = 2^ 6 * ln( 1 +  1 * 2^(- 6+1) + ( 1^2+ 1^2) * 2^(-2* 6) )   n =  6   d_n = 1+1i 
assign u[4'b0101] [07] = 22'h 0001FF;  // +1.9999195675060046 = 2^ 7 * ln( 1 +  1 * 2^(- 7+1) + ( 1^2+ 1^2) * 2^(-2* 7) )   n =  7   d_n = 1+1i 
assign u[4'b0101] [08] = 22'h 0001FF;  // +1.9999797737846823 = 2^ 8 * ln( 1 +  1 * 2^(- 8+1) + ( 1^2+ 1^2) * 2^(-2* 8) )   n =  8   d_n = 1+1i 
assign u[4'b0101] [09] = 22'h 0001FF;  // +1.9999949286148679 = 2^ 9 * ln( 1 +  1 * 2^(- 9+1) + ( 1^2+ 1^2) * 2^(-2* 9) )   n =  9   d_n = 1+1i 
assign u[4'b0101] [10] = 22'h 0001FF;  // +1.9999987302952080 = 2^10 * ln( 1 +  1 * 2^(-10+1) + ( 1^2+ 1^2) * 2^(-2*10) )   n = 10   d_n = 1+1i 
assign u[4'b0101] [11] = 22'h 0001FF;  // +1.9999996823413151 = 2^11 * ln( 1 +  1 * 2^(-11+1) + ( 1^2+ 1^2) * 2^(-2*11) )   n = 11   d_n = 1+1i 
assign u[4'b0101] [12] = 22'h 0001FF;  // +1.9999999205562393 = 2^12 * ln( 1 +  1 * 2^(-12+1) + ( 1^2+ 1^2) * 2^(-2*12) )   n = 12   d_n = 1+1i 
assign u[4'b0101] [13] = 22'h 0001FF;  // +1.9999999801340587 = 2^13 * ln( 1 +  1 * 2^(-13+1) + ( 1^2+ 1^2) * 2^(-2*13) )   n = 13   d_n = 1+1i 
assign u[4'b0101] [14] = 22'h 0001FF;  // +1.9999999950332306 = 2^14 * ln( 1 +  1 * 2^(-14+1) + ( 1^2+ 1^2) * 2^(-2*14) )   n = 14   d_n = 1+1i 
assign u[4'b0101] [15] = 22'h 0001FF;  // +1.9999999987582722 = 2^15 * ln( 1 +  1 * 2^(-15+1) + ( 1^2+ 1^2) * 2^(-2*15) )   n = 15   d_n = 1+1i 
assign u[4'b0101] [16] = 22'h 0001FF;  // +1.9999999996895637 = 2^16 * ln( 1 +  1 * 2^(-16+1) + ( 1^2+ 1^2) * 2^(-2*16) )   n = 16   d_n = 1+1i 
assign u[4'b0101] [17] = 22'h 0001FF;  // +1.9999999999223903 = 2^17 * ln( 1 +  1 * 2^(-17+1) + ( 1^2+ 1^2) * 2^(-2*17) )   n = 17   d_n = 1+1i 
assign u[4'b0101] [18] = 22'h 0001FF;  // +1.9999999999951494 = 2^18 * ln( 1 +  1 * 2^(-18+1) + ( 1^2+ 1^2) * 2^(-2*18) )   n = 18   d_n = 1+1i 
assign u[4'b0101] [19] = 22'h 0001FF;  // +1.9999999999987874 = 2^19 * ln( 1 +  1 * 2^(-19+1) + ( 1^2+ 1^2) * 2^(-2*19) )   n = 19   d_n = 1+1i 
assign u[4'b0101] [20] = 22'h 0001FF;  // +1.9999999999996969 = 2^20 * ln( 1 +  1 * 2^(-20+1) + ( 1^2+ 1^2) * 2^(-2*20) )   n = 20   d_n = 1+1i 
assign u[4'b0101] [21] = 22'h 0001FF;  // +1.9999999999999243 = 2^21 * ln( 1 +  1 * 2^(-21+1) + ( 1^2+ 1^2) * 2^(-2*21) )   n = 21   d_n = 1+1i 
assign u[4'b0101] [22] = 22'h 0001FF;  // +1.9999999999999811 = 2^22 * ln( 1 +  1 * 2^(-22+1) + ( 1^2+ 1^2) * 2^(-2*22) )   n = 22   d_n = 1+1i 
assign u[4'b0101] [23] = 22'h 0001FF;  // +1.9999999999999953 = 2^23 * ln( 1 +  1 * 2^(-23+1) + ( 1^2+ 1^2) * 2^(-2*23) )   n = 23   d_n = 1+1i 
assign u[4'b0101] [24] = 22'h 0001FF;  // +1.9999999999999989 = 2^24 * ln( 1 +  1 * 2^(-24+1) + ( 1^2+ 1^2) * 2^(-2*24) )   n = 24   d_n = 1+1i 
assign u[4'b0101] [25] = 22'h 0001FF;  // +1.9999999999999998 = 2^25 * ln( 1 +  1 * 2^(-25+1) + ( 1^2+ 1^2) * 2^(-2*25) )   n = 25   d_n = 1+1i 
assign u[4'b0101] [26] = 22'h 0001FF;  // +1.9999999850988390 = 2^26 * ln( 1 +  1 * 2^(-26+1) + ( 1^2+ 1^2) * 2^(-2*26) )   n = 26   d_n = 1+1i 
assign u[4'b0101] [27] = 22'h 0001FF;  // +1.9999999925494194 = 2^27 * ln( 1 +  1 * 2^(-27+1) + ( 1^2+ 1^2) * 2^(-2*27) )   n = 27   d_n = 1+1i 
assign u[4'b0101] [28] = 22'h 0001FF;  // +1.9999999962747097 = 2^28 * ln( 1 +  1 * 2^(-28+1) + ( 1^2+ 1^2) * 2^(-2*28) )   n = 28   d_n = 1+1i 
assign u[4'b0101] [29] = 22'h 0001FF;  // +1.9999999981373549 = 2^29 * ln( 1 +  1 * 2^(-29+1) + ( 1^2+ 1^2) * 2^(-2*29) )   n = 29   d_n = 1+1i 
assign u[4'b0101] [30] = 22'h 0001FF;  // +1.9999999990686774 = 2^30 * ln( 1 +  1 * 2^(-30+1) + ( 1^2+ 1^2) * 2^(-2*30) )   n = 30   d_n = 1+1i 
assign u[4'b0101] [31] = 22'h 0001FF;  // +1.9999999995343387 = 2^31 * ln( 1 +  1 * 2^(-31+1) + ( 1^2+ 1^2) * 2^(-2*31) )   n = 31   d_n = 1+1i 
assign u[4'b0101] [32] = 22'h 0001FF;  // +1.9999999997671694 = 2^32 * ln( 1 +  1 * 2^(-32+1) + ( 1^2+ 1^2) * 2^(-2*32) )   n = 32   d_n = 1+1i 
assign u[4'b0101] [33] = 22'h 0001FF;  // +1.9999999998835847 = 2^33 * ln( 1 +  1 * 2^(-33+1) + ( 1^2+ 1^2) * 2^(-2*33) )   n = 33   d_n = 1+1i 
assign u[4'b0101] [34] = 22'h 0001FF;  // +1.9999999999417923 = 2^34 * ln( 1 +  1 * 2^(-34+1) + ( 1^2+ 1^2) * 2^(-2*34) )   n = 34   d_n = 1+1i 
assign u[4'b0101] [35] = 22'h 0001FF;  // +1.9999999999708962 = 2^35 * ln( 1 +  1 * 2^(-35+1) + ( 1^2+ 1^2) * 2^(-2*35) )   n = 35   d_n = 1+1i 
assign u[4'b0101] [36] = 22'h 0001FF;  // +1.9999999999854481 = 2^36 * ln( 1 +  1 * 2^(-36+1) + ( 1^2+ 1^2) * 2^(-2*36) )   n = 36   d_n = 1+1i 
assign u[4'b0101] [37] = 22'h 0001FF;  // +1.9999999999927240 = 2^37 * ln( 1 +  1 * 2^(-37+1) + ( 1^2+ 1^2) * 2^(-2*37) )   n = 37   d_n = 1+1i 
assign u[4'b0101] [38] = 22'h 0001FF;  // +1.9999999999963620 = 2^38 * ln( 1 +  1 * 2^(-38+1) + ( 1^2+ 1^2) * 2^(-2*38) )   n = 38   d_n = 1+1i 
assign u[4'b0101] [39] = 22'h 0001FF;  // +1.9999999999981810 = 2^39 * ln( 1 +  1 * 2^(-39+1) + ( 1^2+ 1^2) * 2^(-2*39) )   n = 39   d_n = 1+1i 
assign u[4'b0101] [40] = 22'h 0001FF;  // +1.9999999999990905 = 2^40 * ln( 1 +  1 * 2^(-40+1) + ( 1^2+ 1^2) * 2^(-2*40) )   n = 40   d_n = 1+1i 
assign u[4'b0101] [41] = 22'h 0001FF;  // +1.9999999999995453 = 2^41 * ln( 1 +  1 * 2^(-41+1) + ( 1^2+ 1^2) * 2^(-2*41) )   n = 41   d_n = 1+1i 
assign u[4'b0101] [42] = 22'h 0001FF;  // +1.9999999999997726 = 2^42 * ln( 1 +  1 * 2^(-42+1) + ( 1^2+ 1^2) * 2^(-2*42) )   n = 42   d_n = 1+1i 
assign u[4'b0101] [43] = 22'h 0001FF;  // +1.9999999999998863 = 2^43 * ln( 1 +  1 * 2^(-43+1) + ( 1^2+ 1^2) * 2^(-2*43) )   n = 43   d_n = 1+1i 
assign u[4'b0101] [44] = 22'h 0001FF;  // +1.9999999999999432 = 2^44 * ln( 1 +  1 * 2^(-44+1) + ( 1^2+ 1^2) * 2^(-2*44) )   n = 44   d_n = 1+1i 
assign u[4'b0101] [45] = 22'h 0001FF;  // +1.9999999999999716 = 2^45 * ln( 1 +  1 * 2^(-45+1) + ( 1^2+ 1^2) * 2^(-2*45) )   n = 45   d_n = 1+1i 
assign u[4'b0101] [46] = 22'h 0001FF;  // +1.9999999999999858 = 2^46 * ln( 1 +  1 * 2^(-46+1) + ( 1^2+ 1^2) * 2^(-2*46) )   n = 46   d_n = 1+1i 
assign u[4'b0101] [47] = 22'h 0001FF;  // +1.9999999999999929 = 2^47 * ln( 1 +  1 * 2^(-47+1) + ( 1^2+ 1^2) * 2^(-2*47) )   n = 47   d_n = 1+1i 
assign u[4'b0101] [48] = 22'h 0001FF;  // +1.9999999999999964 = 2^48 * ln( 1 +  1 * 2^(-48+1) + ( 1^2+ 1^2) * 2^(-2*48) )   n = 48   d_n = 1+1i 
assign u[4'b0101] [49] = 22'h 0001FF;  // +1.9999999999999982 = 2^49 * ln( 1 +  1 * 2^(-49+1) + ( 1^2+ 1^2) * 2^(-2*49) )   n = 49   d_n = 1+1i 
assign u[4'b0101] [50] = 22'h 0001FF;  // +1.9999999999999991 = 2^50 * ln( 1 +  1 * 2^(-50+1) + ( 1^2+ 1^2) * 2^(-2*50) )   n = 50   d_n = 1+1i 
assign u[4'b0101] [51] = 22'h 0001FF;  // +1.9999999999999996 = 2^51 * ln( 1 +  1 * 2^(-51+1) + ( 1^2+ 1^2) * 2^(-2*51) )   n = 51   d_n = 1+1i 
assign u[4'b0101] [52] = 22'h 0001FF;  // +1.9999999999999998 = 2^52 * ln( 1 +  1 * 2^(-52+1) + ( 1^2+ 1^2) * 2^(-2*52) )   n = 52   d_n = 1+1i 
assign u[4'b0101] [53] = 22'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  1 * 2^(-53+1) + ( 1^2+ 1^2) * 2^(-2*53) )   n = 53   d_n = 1+1i 
assign u[4'b0101] [54] = 22'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  1 * 2^(-54+1) + ( 1^2+ 1^2) * 2^(-2*54) )   n = 54   d_n = 1+1i 
assign u[4'b0101] [55] = 22'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  1 * 2^(-55+1) + ( 1^2+ 1^2) * 2^(-2*55) )   n = 55   d_n = 1+1i 
assign u[4'b0101] [56] = 22'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  1 * 2^(-56+1) + ( 1^2+ 1^2) * 2^(-2*56) )   n = 56   d_n = 1+1i 
assign u[4'b0101] [57] = 22'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  1 * 2^(-57+1) + ( 1^2+ 1^2) * 2^(-2*57) )   n = 57   d_n = 1+1i 
assign u[4'b0101] [58] = 22'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  1 * 2^(-58+1) + ( 1^2+ 1^2) * 2^(-2*58) )   n = 58   d_n = 1+1i 
assign u[4'b0101] [59] = 22'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  1 * 2^(-59+1) + ( 1^2+ 1^2) * 2^(-2*59) )   n = 59   d_n = 1+1i 
assign u[4'b0101] [60] = 22'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  1 * 2^(-60+1) + ( 1^2+ 1^2) * 2^(-2*60) )   n = 60   d_n = 1+1i 
assign u[4'b0101] [61] = 22'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  1 * 2^(-61+1) + ( 1^2+ 1^2) * 2^(-2*61) )   n = 61   d_n = 1+1i 
assign u[4'b0101] [62] = 22'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  1 * 2^(-62+1) + ( 1^2+ 1^2) * 2^(-2*62) )   n = 62   d_n = 1+1i 
assign u[4'b0101] [63] = 22'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  1 * 2^(-63+1) + ( 1^2+ 1^2) * 2^(-2*63) )   n = 63   d_n = 1+1i 
assign u[4'b0101] [64] = 22'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  1 * 2^(-64+1) + ( 1^2+ 1^2) * 2^(-2*64) )   n = 64   d_n = 1+1i 
assign u[4'b0110] [01] = 22'h 000072;  // +0.4462871026284197 = 2^ 1 * ln( 1 +  0 * 2^(- 1+1) + ( 0^2+ 1^2) * 2^(-2* 1) )   n =  1   d_n = 0+1i 
assign u[4'b0110] [02] = 22'h 00003E;  // +0.2424984872657394 = 2^ 2 * ln( 1 +  0 * 2^(- 2+1) + ( 0^2+ 1^2) * 2^(-2* 2) )   n =  2   d_n = 0+1i 
assign u[4'b0110] [03] = 22'h 00001F;  // +0.1240334922877210 = 2^ 3 * ln( 1 +  0 * 2^(- 3+1) + ( 0^2+ 1^2) * 2^(-2* 3) )   n =  3   d_n = 0+1i 
assign u[4'b0110] [04] = 22'h 00000F;  // +0.0623782466505195 = 2^ 4 * ln( 1 +  0 * 2^(- 4+1) + ( 0^2+ 1^2) * 2^(-2* 4) )   n =  4   d_n = 0+1i 
assign u[4'b0110] [05] = 22'h 000007;  // +0.0312347511377731 = 2^ 5 * ln( 1 +  0 * 2^(- 5+1) + ( 0^2+ 1^2) * 2^(-2* 5) )   n =  5   d_n = 0+1i 
assign u[4'b0110] [06] = 22'h 000003;  // +0.0156230929617406 = 2^ 6 * ln( 1 +  0 * 2^(- 6+1) + ( 0^2+ 1^2) * 2^(-2* 6) )   n =  6   d_n = 0+1i 
assign u[4'b0110] [07] = 22'h 000001;  // +0.0078122615911219 = 2^ 7 * ln( 1 +  0 * 2^(- 7+1) + ( 0^2+ 1^2) * 2^(-2* 7) )   n =  7   d_n = 0+1i 
assign u[4'b0110] [08] = 22'h 000000;  // +0.0039062201979808 = 2^ 8 * ln( 1 +  0 * 2^(- 8+1) + ( 0^2+ 1^2) * 2^(-2* 8) )   n =  8   d_n = 0+1i 
assign u[4'b0110] [09] = 22'h 000000;  // +0.0019531212747156 = 2^ 9 * ln( 1 +  0 * 2^(- 9+1) + ( 0^2+ 1^2) * 2^(-2* 9) )   n =  9   d_n = 0+1i 
assign u[4'b0110] [10] = 22'h 000000;  // +0.0009765620343389 = 2^10 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 1^2) * 2^(-2*10) )   n = 10   d_n = 0+1i 
assign u[4'b0110] [11] = 22'h 000000;  // +0.0004882811917923 = 2^11 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 1^2) * 2^(-2*11) )   n = 11   d_n = 0+1i 
assign u[4'b0110] [12] = 22'h 000000;  // +0.0002441406177240 = 2^12 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 1^2) * 2^(-2*12) )   n = 12   d_n = 0+1i 
assign u[4'b0110] [13] = 22'h 000000;  // +0.0001220703120453 = 2^13 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 1^2) * 2^(-2*13) )   n = 13   d_n = 0+1i 
assign u[4'b0110] [14] = 22'h 000000;  // +0.0000610351561932 = 2^14 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 1^2) * 2^(-2*14) )   n = 14   d_n = 0+1i 
assign u[4'b0110] [15] = 22'h 000000;  // +0.0000305175781179 = 2^15 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 1^2) * 2^(-2*15) )   n = 15   d_n = 0+1i 
assign u[4'b0110] [16] = 22'h 000000;  // +0.0000152587890616 = 2^16 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 1^2) * 2^(-2*16) )   n = 16   d_n = 0+1i 
assign u[4'b0110] [17] = 22'h 000000;  // +0.0000076293945311 = 2^17 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 1^2) * 2^(-2*17) )   n = 17   d_n = 0+1i 
assign u[4'b0110] [18] = 22'h 000000;  // +0.0000038146972656 = 2^18 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 1^2) * 2^(-2*18) )   n = 18   d_n = 0+1i 
assign u[4'b0110] [19] = 22'h 000000;  // +0.0000019073486328 = 2^19 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 1^2) * 2^(-2*19) )   n = 19   d_n = 0+1i 
assign u[4'b0110] [20] = 22'h 000000;  // +0.0000009536743164 = 2^20 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 1^2) * 2^(-2*20) )   n = 20   d_n = 0+1i 
assign u[4'b0110] [21] = 22'h 000000;  // +0.0000004768371582 = 2^21 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 1^2) * 2^(-2*21) )   n = 21   d_n = 0+1i 
assign u[4'b0110] [22] = 22'h 000000;  // +0.0000002384185791 = 2^22 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 1^2) * 2^(-2*22) )   n = 22   d_n = 0+1i 
assign u[4'b0110] [23] = 22'h 000000;  // +0.0000001192092896 = 2^23 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 1^2) * 2^(-2*23) )   n = 23   d_n = 0+1i 
assign u[4'b0110] [24] = 22'h 000000;  // +0.0000000596046448 = 2^24 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 1^2) * 2^(-2*24) )   n = 24   d_n = 0+1i 
assign u[4'b0110] [25] = 22'h 000000;  // +0.0000000298023224 = 2^25 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 1^2) * 2^(-2*25) )   n = 25   d_n = 0+1i 
assign u[4'b0110] [26] = 22'h 000000;  // +0.0000000000000000 = 2^26 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 1^2) * 2^(-2*26) )   n = 26   d_n = 0+1i 
assign u[4'b0110] [27] = 22'h 000000;  // +0.0000000000000000 = 2^27 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 1^2) * 2^(-2*27) )   n = 27   d_n = 0+1i 
assign u[4'b0110] [28] = 22'h 000000;  // +0.0000000000000000 = 2^28 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 1^2) * 2^(-2*28) )   n = 28   d_n = 0+1i 
assign u[4'b0110] [29] = 22'h 000000;  // +0.0000000000000000 = 2^29 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 1^2) * 2^(-2*29) )   n = 29   d_n = 0+1i 
assign u[4'b0110] [30] = 22'h 000000;  // +0.0000000000000000 = 2^30 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 1^2) * 2^(-2*30) )   n = 30   d_n = 0+1i 
assign u[4'b0110] [31] = 22'h 000000;  // +0.0000000000000000 = 2^31 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 1^2) * 2^(-2*31) )   n = 31   d_n = 0+1i 
assign u[4'b0110] [32] = 22'h 000000;  // +0.0000000000000000 = 2^32 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 1^2) * 2^(-2*32) )   n = 32   d_n = 0+1i 
assign u[4'b0110] [33] = 22'h 000000;  // +0.0000000000000000 = 2^33 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 1^2) * 2^(-2*33) )   n = 33   d_n = 0+1i 
assign u[4'b0110] [34] = 22'h 000000;  // +0.0000000000000000 = 2^34 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 1^2) * 2^(-2*34) )   n = 34   d_n = 0+1i 
assign u[4'b0110] [35] = 22'h 000000;  // +0.0000000000000000 = 2^35 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 1^2) * 2^(-2*35) )   n = 35   d_n = 0+1i 
assign u[4'b0110] [36] = 22'h 000000;  // +0.0000000000000000 = 2^36 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 1^2) * 2^(-2*36) )   n = 36   d_n = 0+1i 
assign u[4'b0110] [37] = 22'h 000000;  // +0.0000000000000000 = 2^37 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 1^2) * 2^(-2*37) )   n = 37   d_n = 0+1i 
assign u[4'b0110] [38] = 22'h 000000;  // +0.0000000000000000 = 2^38 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 1^2) * 2^(-2*38) )   n = 38   d_n = 0+1i 
assign u[4'b0110] [39] = 22'h 000000;  // +0.0000000000000000 = 2^39 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 1^2) * 2^(-2*39) )   n = 39   d_n = 0+1i 
assign u[4'b0110] [40] = 22'h 000000;  // +0.0000000000000000 = 2^40 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 1^2) * 2^(-2*40) )   n = 40   d_n = 0+1i 
assign u[4'b0110] [41] = 22'h 000000;  // +0.0000000000000000 = 2^41 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 1^2) * 2^(-2*41) )   n = 41   d_n = 0+1i 
assign u[4'b0110] [42] = 22'h 000000;  // +0.0000000000000000 = 2^42 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 1^2) * 2^(-2*42) )   n = 42   d_n = 0+1i 
assign u[4'b0110] [43] = 22'h 000000;  // +0.0000000000000000 = 2^43 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 1^2) * 2^(-2*43) )   n = 43   d_n = 0+1i 
assign u[4'b0110] [44] = 22'h 000000;  // +0.0000000000000000 = 2^44 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 1^2) * 2^(-2*44) )   n = 44   d_n = 0+1i 
assign u[4'b0110] [45] = 22'h 000000;  // +0.0000000000000000 = 2^45 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 1^2) * 2^(-2*45) )   n = 45   d_n = 0+1i 
assign u[4'b0110] [46] = 22'h 000000;  // +0.0000000000000000 = 2^46 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 1^2) * 2^(-2*46) )   n = 46   d_n = 0+1i 
assign u[4'b0110] [47] = 22'h 000000;  // +0.0000000000000000 = 2^47 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 1^2) * 2^(-2*47) )   n = 47   d_n = 0+1i 
assign u[4'b0110] [48] = 22'h 000000;  // +0.0000000000000000 = 2^48 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 1^2) * 2^(-2*48) )   n = 48   d_n = 0+1i 
assign u[4'b0110] [49] = 22'h 000000;  // +0.0000000000000000 = 2^49 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 1^2) * 2^(-2*49) )   n = 49   d_n = 0+1i 
assign u[4'b0110] [50] = 22'h 000000;  // +0.0000000000000000 = 2^50 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 1^2) * 2^(-2*50) )   n = 50   d_n = 0+1i 
assign u[4'b0110] [51] = 22'h 000000;  // +0.0000000000000000 = 2^51 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 1^2) * 2^(-2*51) )   n = 51   d_n = 0+1i 
assign u[4'b0110] [52] = 22'h 000000;  // +0.0000000000000000 = 2^52 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 1^2) * 2^(-2*52) )   n = 52   d_n = 0+1i 
assign u[4'b0110] [53] = 22'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 1^2) * 2^(-2*53) )   n = 53   d_n = 0+1i 
assign u[4'b0110] [54] = 22'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 1^2) * 2^(-2*54) )   n = 54   d_n = 0+1i 
assign u[4'b0110] [55] = 22'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 1^2) * 2^(-2*55) )   n = 55   d_n = 0+1i 
assign u[4'b0110] [56] = 22'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 1^2) * 2^(-2*56) )   n = 56   d_n = 0+1i 
assign u[4'b0110] [57] = 22'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 1^2) * 2^(-2*57) )   n = 57   d_n = 0+1i 
assign u[4'b0110] [58] = 22'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 1^2) * 2^(-2*58) )   n = 58   d_n = 0+1i 
assign u[4'b0110] [59] = 22'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 1^2) * 2^(-2*59) )   n = 59   d_n = 0+1i 
assign u[4'b0110] [60] = 22'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 1^2) * 2^(-2*60) )   n = 60   d_n = 0+1i 
assign u[4'b0110] [61] = 22'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 1^2) * 2^(-2*61) )   n = 61   d_n = 0+1i 
assign u[4'b0110] [62] = 22'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 1^2) * 2^(-2*62) )   n = 62   d_n = 0+1i 
assign u[4'b0110] [63] = 22'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 1^2) * 2^(-2*63) )   n = 63   d_n = 0+1i 
assign u[4'b0110] [64] = 22'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 1^2) * 2^(-2*64) )   n = 64   d_n = 0+1i 
assign u[4'b0111] [01] = 22'h 3FFE9D;  // -1.3862943611198904 = 2^ 1 * ln( 1 + -1 * 2^(- 1+1) + (-1^2+ 1^2) * 2^(-2* 1) )   n =  1   d_n = -1+1i 
assign u[4'b0111] [02] = 22'h 3FFE1E;  // -1.8800145169829416 = 2^ 2 * ln( 1 + -1 * 2^(- 2+1) + (-1^2+ 1^2) * 2^(-2* 2) )   n =  2   d_n = -1+1i 
assign u[4'b0111] [03] = 22'h 3FFE06;  // -1.9748806234522058 = 2^ 3 * ln( 1 + -1 * 2^(- 3+1) + (-1^2+ 1^2) * 2^(-2* 3) )   n =  3   d_n = -1+1i 
assign u[4'b0111] [04] = 22'h 3FFE01;  // -1.9942791233164259 = 2^ 4 * ln( 1 + -1 * 2^(- 4+1) + (-1^2+ 1^2) * 2^(-2* 4) )   n =  4   d_n = -1+1i 
assign u[4'b0111] [05] = 22'h 3FFE00;  // -1.9986353578798890 = 2^ 5 * ln( 1 + -1 * 2^(- 5+1) + (-1^2+ 1^2) * 2^(-2* 5) )   n =  5   d_n = -1+1i 
assign u[4'b0111] [06] = 22'h 3FFE00;  // -1.9996667544388824 = 2^ 6 * ln( 1 + -1 * 2^(- 6+1) + (-1^2+ 1^2) * 2^(-2* 6) )   n =  6   d_n = -1+1i 
assign u[4'b0111] [07] = 22'h 3FFE00;  // -1.9999176601574109 = 2^ 7 * ln( 1 + -1 * 2^(- 7+1) + (-1^2+ 1^2) * 2^(-2* 7) )   n =  7   d_n = -1+1i 
assign u[4'b0111] [08] = 22'h 3FFE00;  // -1.9999795353661032 = 2^ 8 * ln( 1 + -1 * 2^(- 8+1) + (-1^2+ 1^2) * 2^(-2* 8) )   n =  8   d_n = -1+1i 
assign u[4'b0111] [09] = 22'h 3FFE00;  // -1.9999948988125242 = 2^ 9 * ln( 1 + -1 * 2^(- 9+1) + (-1^2+ 1^2) * 2^(-2* 9) )   n =  9   d_n = -1+1i 
assign u[4'b0111] [10] = 22'h 3FFE00;  // -1.9999987265701442 = 2^10 * ln( 1 + -1 * 2^(-10+1) + (-1^2+ 1^2) * 2^(-2*10) )   n = 10   d_n = -1+1i 
assign u[4'b0111] [11] = 22'h 3FFE00;  // -1.9999996818756538 = 2^11 * ln( 1 + -1 * 2^(-11+1) + (-1^2+ 1^2) * 2^(-2*11) )   n = 11   d_n = -1+1i 
assign u[4'b0111] [12] = 22'h 3FFE00;  // -1.9999999204980317 = 2^12 * ln( 1 + -1 * 2^(-12+1) + (-1^2+ 1^2) * 2^(-2*12) )   n = 12   d_n = -1+1i 
assign u[4'b0111] [13] = 22'h 3FFE00;  // -1.9999999801276920 = 2^13 * ln( 1 + -1 * 2^(-13+1) + (-1^2+ 1^2) * 2^(-2*13) )   n = 13   d_n = -1+1i 
assign u[4'b0111] [14] = 22'h 3FFE00;  // -1.9999999950326621 = 2^14 * ln( 1 + -1 * 2^(-14+1) + (-1^2+ 1^2) * 2^(-2*14) )   n = 14   d_n = -1+1i 
assign u[4'b0111] [15] = 22'h 3FFE00;  // -1.9999999987582011 = 2^15 * ln( 1 + -1 * 2^(-15+1) + (-1^2+ 1^2) * 2^(-2*15) )   n = 15   d_n = -1+1i 
assign u[4'b0111] [16] = 22'h 3FFE00;  // -1.9999999996895548 = 2^16 * ln( 1 + -1 * 2^(-16+1) + (-1^2+ 1^2) * 2^(-2*16) )   n = 16   d_n = -1+1i 
assign u[4'b0111] [17] = 22'h 3FFE00;  // -1.9999999999223892 = 2^17 * ln( 1 + -1 * 2^(-17+1) + (-1^2+ 1^2) * 2^(-2*17) )   n = 17   d_n = -1+1i 
assign u[4'b0111] [18] = 22'h 3FFE00;  // -1.9999999999951494 = 2^18 * ln( 1 + -1 * 2^(-18+1) + (-1^2+ 1^2) * 2^(-2*18) )   n = 18   d_n = -1+1i 
assign u[4'b0111] [19] = 22'h 3FFE00;  // -1.9999999999987874 = 2^19 * ln( 1 + -1 * 2^(-19+1) + (-1^2+ 1^2) * 2^(-2*19) )   n = 19   d_n = -1+1i 
assign u[4'b0111] [20] = 22'h 3FFE00;  // -1.9999999999996969 = 2^20 * ln( 1 + -1 * 2^(-20+1) + (-1^2+ 1^2) * 2^(-2*20) )   n = 20   d_n = -1+1i 
assign u[4'b0111] [21] = 22'h 3FFE00;  // -1.9999999999999243 = 2^21 * ln( 1 + -1 * 2^(-21+1) + (-1^2+ 1^2) * 2^(-2*21) )   n = 21   d_n = -1+1i 
assign u[4'b0111] [22] = 22'h 3FFE00;  // -1.9999999999999811 = 2^22 * ln( 1 + -1 * 2^(-22+1) + (-1^2+ 1^2) * 2^(-2*22) )   n = 22   d_n = -1+1i 
assign u[4'b0111] [23] = 22'h 3FFE00;  // -1.9999999999999953 = 2^23 * ln( 1 + -1 * 2^(-23+1) + (-1^2+ 1^2) * 2^(-2*23) )   n = 23   d_n = -1+1i 
assign u[4'b0111] [24] = 22'h 3FFE00;  // -1.9999999999999989 = 2^24 * ln( 1 + -1 * 2^(-24+1) + (-1^2+ 1^2) * 2^(-2*24) )   n = 24   d_n = -1+1i 
assign u[4'b0111] [25] = 22'h 3FFE00;  // -1.9999999999999998 = 2^25 * ln( 1 + -1 * 2^(-25+1) + (-1^2+ 1^2) * 2^(-2*25) )   n = 25   d_n = -1+1i 
assign u[4'b0111] [26] = 22'h 3FFE00;  // -2.0000000000000000 = 2^26 * ln( 1 + -1 * 2^(-26+1) + (-1^2+ 1^2) * 2^(-2*26) )   n = 26   d_n = -1+1i 
assign u[4'b0111] [27] = 22'h 3FFDFF;  // -2.0000000074505806 = 2^27 * ln( 1 + -1 * 2^(-27+1) + (-1^2+ 1^2) * 2^(-2*27) )   n = 27   d_n = -1+1i 
assign u[4'b0111] [28] = 22'h 3FFDFF;  // -2.0000000037252903 = 2^28 * ln( 1 + -1 * 2^(-28+1) + (-1^2+ 1^2) * 2^(-2*28) )   n = 28   d_n = -1+1i 
assign u[4'b0111] [29] = 22'h 3FFDFF;  // -2.0000000018626451 = 2^29 * ln( 1 + -1 * 2^(-29+1) + (-1^2+ 1^2) * 2^(-2*29) )   n = 29   d_n = -1+1i 
assign u[4'b0111] [30] = 22'h 3FFDFF;  // -2.0000000009313226 = 2^30 * ln( 1 + -1 * 2^(-30+1) + (-1^2+ 1^2) * 2^(-2*30) )   n = 30   d_n = -1+1i 
assign u[4'b0111] [31] = 22'h 3FFDFF;  // -2.0000000004656613 = 2^31 * ln( 1 + -1 * 2^(-31+1) + (-1^2+ 1^2) * 2^(-2*31) )   n = 31   d_n = -1+1i 
assign u[4'b0111] [32] = 22'h 3FFDFF;  // -2.0000000002328306 = 2^32 * ln( 1 + -1 * 2^(-32+1) + (-1^2+ 1^2) * 2^(-2*32) )   n = 32   d_n = -1+1i 
assign u[4'b0111] [33] = 22'h 3FFDFF;  // -2.0000000001164153 = 2^33 * ln( 1 + -1 * 2^(-33+1) + (-1^2+ 1^2) * 2^(-2*33) )   n = 33   d_n = -1+1i 
assign u[4'b0111] [34] = 22'h 3FFDFF;  // -2.0000000000582077 = 2^34 * ln( 1 + -1 * 2^(-34+1) + (-1^2+ 1^2) * 2^(-2*34) )   n = 34   d_n = -1+1i 
assign u[4'b0111] [35] = 22'h 3FFDFF;  // -2.0000000000291038 = 2^35 * ln( 1 + -1 * 2^(-35+1) + (-1^2+ 1^2) * 2^(-2*35) )   n = 35   d_n = -1+1i 
assign u[4'b0111] [36] = 22'h 3FFDFF;  // -2.0000000000145519 = 2^36 * ln( 1 + -1 * 2^(-36+1) + (-1^2+ 1^2) * 2^(-2*36) )   n = 36   d_n = -1+1i 
assign u[4'b0111] [37] = 22'h 3FFDFF;  // -2.0000000000072760 = 2^37 * ln( 1 + -1 * 2^(-37+1) + (-1^2+ 1^2) * 2^(-2*37) )   n = 37   d_n = -1+1i 
assign u[4'b0111] [38] = 22'h 3FFDFF;  // -2.0000000000036380 = 2^38 * ln( 1 + -1 * 2^(-38+1) + (-1^2+ 1^2) * 2^(-2*38) )   n = 38   d_n = -1+1i 
assign u[4'b0111] [39] = 22'h 3FFDFF;  // -2.0000000000018190 = 2^39 * ln( 1 + -1 * 2^(-39+1) + (-1^2+ 1^2) * 2^(-2*39) )   n = 39   d_n = -1+1i 
assign u[4'b0111] [40] = 22'h 3FFE00;  // -2.0000000000009095 = 2^40 * ln( 1 + -1 * 2^(-40+1) + (-1^2+ 1^2) * 2^(-2*40) )   n = 40   d_n = -1+1i 
assign u[4'b0111] [41] = 22'h 3FFE00;  // -2.0000000000004547 = 2^41 * ln( 1 + -1 * 2^(-41+1) + (-1^2+ 1^2) * 2^(-2*41) )   n = 41   d_n = -1+1i 
assign u[4'b0111] [42] = 22'h 3FFE00;  // -2.0000000000002274 = 2^42 * ln( 1 + -1 * 2^(-42+1) + (-1^2+ 1^2) * 2^(-2*42) )   n = 42   d_n = -1+1i 
assign u[4'b0111] [43] = 22'h 3FFE00;  // -2.0000000000001137 = 2^43 * ln( 1 + -1 * 2^(-43+1) + (-1^2+ 1^2) * 2^(-2*43) )   n = 43   d_n = -1+1i 
assign u[4'b0111] [44] = 22'h 3FFE00;  // -2.0000000000000568 = 2^44 * ln( 1 + -1 * 2^(-44+1) + (-1^2+ 1^2) * 2^(-2*44) )   n = 44   d_n = -1+1i 
assign u[4'b0111] [45] = 22'h 3FFE00;  // -2.0000000000000284 = 2^45 * ln( 1 + -1 * 2^(-45+1) + (-1^2+ 1^2) * 2^(-2*45) )   n = 45   d_n = -1+1i 
assign u[4'b0111] [46] = 22'h 3FFE00;  // -2.0000000000000142 = 2^46 * ln( 1 + -1 * 2^(-46+1) + (-1^2+ 1^2) * 2^(-2*46) )   n = 46   d_n = -1+1i 
assign u[4'b0111] [47] = 22'h 3FFE00;  // -2.0000000000000071 = 2^47 * ln( 1 + -1 * 2^(-47+1) + (-1^2+ 1^2) * 2^(-2*47) )   n = 47   d_n = -1+1i 
assign u[4'b0111] [48] = 22'h 3FFE00;  // -2.0000000000000036 = 2^48 * ln( 1 + -1 * 2^(-48+1) + (-1^2+ 1^2) * 2^(-2*48) )   n = 48   d_n = -1+1i 
assign u[4'b0111] [49] = 22'h 3FFE00;  // -2.0000000000000018 = 2^49 * ln( 1 + -1 * 2^(-49+1) + (-1^2+ 1^2) * 2^(-2*49) )   n = 49   d_n = -1+1i 
assign u[4'b0111] [50] = 22'h 3FFE00;  // -2.0000000000000009 = 2^50 * ln( 1 + -1 * 2^(-50+1) + (-1^2+ 1^2) * 2^(-2*50) )   n = 50   d_n = -1+1i 
assign u[4'b0111] [51] = 22'h 3FFE00;  // -2.0000000000000004 = 2^51 * ln( 1 + -1 * 2^(-51+1) + (-1^2+ 1^2) * 2^(-2*51) )   n = 51   d_n = -1+1i 
assign u[4'b0111] [52] = 22'h 3FFE00;  // -2.0000000000000004 = 2^52 * ln( 1 + -1 * 2^(-52+1) + (-1^2+ 1^2) * 2^(-2*52) )   n = 52   d_n = -1+1i 
assign u[4'b0111] [53] = 22'h 3FFE00;  // -2.0000000000000000 = 2^53 * ln( 1 + -1 * 2^(-53+1) + (-1^2+ 1^2) * 2^(-2*53) )   n = 53   d_n = -1+1i 
assign u[4'b0111] [54] = 22'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 + -1 * 2^(-54+1) + (-1^2+ 1^2) * 2^(-2*54) )   n = 54   d_n = -1+1i 
assign u[4'b0111] [55] = 22'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 + -1 * 2^(-55+1) + (-1^2+ 1^2) * 2^(-2*55) )   n = 55   d_n = -1+1i 
assign u[4'b0111] [56] = 22'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 + -1 * 2^(-56+1) + (-1^2+ 1^2) * 2^(-2*56) )   n = 56   d_n = -1+1i 
assign u[4'b0111] [57] = 22'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 + -1 * 2^(-57+1) + (-1^2+ 1^2) * 2^(-2*57) )   n = 57   d_n = -1+1i 
assign u[4'b0111] [58] = 22'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 + -1 * 2^(-58+1) + (-1^2+ 1^2) * 2^(-2*58) )   n = 58   d_n = -1+1i 
assign u[4'b0111] [59] = 22'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 + -1 * 2^(-59+1) + (-1^2+ 1^2) * 2^(-2*59) )   n = 59   d_n = -1+1i 
assign u[4'b0111] [60] = 22'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 + -1 * 2^(-60+1) + (-1^2+ 1^2) * 2^(-2*60) )   n = 60   d_n = -1+1i 
assign u[4'b0111] [61] = 22'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 + -1 * 2^(-61+1) + (-1^2+ 1^2) * 2^(-2*61) )   n = 61   d_n = -1+1i 
assign u[4'b0111] [62] = 22'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 + -1 * 2^(-62+1) + (-1^2+ 1^2) * 2^(-2*62) )   n = 62   d_n = -1+1i 
assign u[4'b0111] [63] = 22'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 + -1 * 2^(-63+1) + (-1^2+ 1^2) * 2^(-2*63) )   n = 63   d_n = -1+1i 
assign u[4'b0111] [64] = 22'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 + -1 * 2^(-64+1) + (-1^2+ 1^2) * 2^(-2*64) )   n = 64   d_n = -1+1i 
assign u[4'b1000] [01] = 22'h 000000;  // +0.0000000000000000 = 2^ 1 * ln( 1 +  0 * 2^(- 1+1) + ( 0^2+ 0^2) * 2^(-2* 1) )   n =  1   d_n = 0 
assign u[4'b1000] [02] = 22'h 000000;  // +0.0000000000000000 = 2^ 2 * ln( 1 +  0 * 2^(- 2+1) + ( 0^2+ 0^2) * 2^(-2* 2) )   n =  2   d_n = 0 
assign u[4'b1000] [03] = 22'h 000000;  // +0.0000000000000000 = 2^ 3 * ln( 1 +  0 * 2^(- 3+1) + ( 0^2+ 0^2) * 2^(-2* 3) )   n =  3   d_n = 0 
assign u[4'b1000] [04] = 22'h 000000;  // +0.0000000000000000 = 2^ 4 * ln( 1 +  0 * 2^(- 4+1) + ( 0^2+ 0^2) * 2^(-2* 4) )   n =  4   d_n = 0 
assign u[4'b1000] [05] = 22'h 000000;  // +0.0000000000000000 = 2^ 5 * ln( 1 +  0 * 2^(- 5+1) + ( 0^2+ 0^2) * 2^(-2* 5) )   n =  5   d_n = 0 
assign u[4'b1000] [06] = 22'h 000000;  // +0.0000000000000000 = 2^ 6 * ln( 1 +  0 * 2^(- 6+1) + ( 0^2+ 0^2) * 2^(-2* 6) )   n =  6   d_n = 0 
assign u[4'b1000] [07] = 22'h 000000;  // +0.0000000000000000 = 2^ 7 * ln( 1 +  0 * 2^(- 7+1) + ( 0^2+ 0^2) * 2^(-2* 7) )   n =  7   d_n = 0 
assign u[4'b1000] [08] = 22'h 000000;  // +0.0000000000000000 = 2^ 8 * ln( 1 +  0 * 2^(- 8+1) + ( 0^2+ 0^2) * 2^(-2* 8) )   n =  8   d_n = 0 
assign u[4'b1000] [09] = 22'h 000000;  // +0.0000000000000000 = 2^ 9 * ln( 1 +  0 * 2^(- 9+1) + ( 0^2+ 0^2) * 2^(-2* 9) )   n =  9   d_n = 0 
assign u[4'b1000] [10] = 22'h 000000;  // +0.0000000000000000 = 2^10 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = 0 
assign u[4'b1000] [11] = 22'h 000000;  // +0.0000000000000000 = 2^11 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = 0 
assign u[4'b1000] [12] = 22'h 000000;  // +0.0000000000000000 = 2^12 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = 0 
assign u[4'b1000] [13] = 22'h 000000;  // +0.0000000000000000 = 2^13 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = 0 
assign u[4'b1000] [14] = 22'h 000000;  // +0.0000000000000000 = 2^14 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = 0 
assign u[4'b1000] [15] = 22'h 000000;  // +0.0000000000000000 = 2^15 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = 0 
assign u[4'b1000] [16] = 22'h 000000;  // +0.0000000000000000 = 2^16 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = 0 
assign u[4'b1000] [17] = 22'h 000000;  // +0.0000000000000000 = 2^17 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = 0 
assign u[4'b1000] [18] = 22'h 000000;  // +0.0000000000000000 = 2^18 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = 0 
assign u[4'b1000] [19] = 22'h 000000;  // +0.0000000000000000 = 2^19 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = 0 
assign u[4'b1000] [20] = 22'h 000000;  // +0.0000000000000000 = 2^20 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = 0 
assign u[4'b1000] [21] = 22'h 000000;  // +0.0000000000000000 = 2^21 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = 0 
assign u[4'b1000] [22] = 22'h 000000;  // +0.0000000000000000 = 2^22 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = 0 
assign u[4'b1000] [23] = 22'h 000000;  // +0.0000000000000000 = 2^23 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = 0 
assign u[4'b1000] [24] = 22'h 000000;  // +0.0000000000000000 = 2^24 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = 0 
assign u[4'b1000] [25] = 22'h 000000;  // +0.0000000000000000 = 2^25 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = 0 
assign u[4'b1000] [26] = 22'h 000000;  // +0.0000000000000000 = 2^26 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = 0 
assign u[4'b1000] [27] = 22'h 000000;  // +0.0000000000000000 = 2^27 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = 0 
assign u[4'b1000] [28] = 22'h 000000;  // +0.0000000000000000 = 2^28 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = 0 
assign u[4'b1000] [29] = 22'h 000000;  // +0.0000000000000000 = 2^29 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = 0 
assign u[4'b1000] [30] = 22'h 000000;  // +0.0000000000000000 = 2^30 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = 0 
assign u[4'b1000] [31] = 22'h 000000;  // +0.0000000000000000 = 2^31 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = 0 
assign u[4'b1000] [32] = 22'h 000000;  // +0.0000000000000000 = 2^32 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = 0 
assign u[4'b1000] [33] = 22'h 000000;  // +0.0000000000000000 = 2^33 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = 0 
assign u[4'b1000] [34] = 22'h 000000;  // +0.0000000000000000 = 2^34 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = 0 
assign u[4'b1000] [35] = 22'h 000000;  // +0.0000000000000000 = 2^35 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = 0 
assign u[4'b1000] [36] = 22'h 000000;  // +0.0000000000000000 = 2^36 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = 0 
assign u[4'b1000] [37] = 22'h 000000;  // +0.0000000000000000 = 2^37 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = 0 
assign u[4'b1000] [38] = 22'h 000000;  // +0.0000000000000000 = 2^38 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = 0 
assign u[4'b1000] [39] = 22'h 000000;  // +0.0000000000000000 = 2^39 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = 0 
assign u[4'b1000] [40] = 22'h 000000;  // +0.0000000000000000 = 2^40 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = 0 
assign u[4'b1000] [41] = 22'h 000000;  // +0.0000000000000000 = 2^41 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = 0 
assign u[4'b1000] [42] = 22'h 000000;  // +0.0000000000000000 = 2^42 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = 0 
assign u[4'b1000] [43] = 22'h 000000;  // +0.0000000000000000 = 2^43 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = 0 
assign u[4'b1000] [44] = 22'h 000000;  // +0.0000000000000000 = 2^44 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = 0 
assign u[4'b1000] [45] = 22'h 000000;  // +0.0000000000000000 = 2^45 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = 0 
assign u[4'b1000] [46] = 22'h 000000;  // +0.0000000000000000 = 2^46 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = 0 
assign u[4'b1000] [47] = 22'h 000000;  // +0.0000000000000000 = 2^47 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = 0 
assign u[4'b1000] [48] = 22'h 000000;  // +0.0000000000000000 = 2^48 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = 0 
assign u[4'b1000] [49] = 22'h 000000;  // +0.0000000000000000 = 2^49 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = 0 
assign u[4'b1000] [50] = 22'h 000000;  // +0.0000000000000000 = 2^50 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = 0 
assign u[4'b1000] [51] = 22'h 000000;  // +0.0000000000000000 = 2^51 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = 0 
assign u[4'b1000] [52] = 22'h 000000;  // +0.0000000000000000 = 2^52 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = 0 
assign u[4'b1000] [53] = 22'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = 0 
assign u[4'b1000] [54] = 22'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = 0 
assign u[4'b1000] [55] = 22'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = 0 
assign u[4'b1000] [56] = 22'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = 0 
assign u[4'b1000] [57] = 22'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = 0 
assign u[4'b1000] [58] = 22'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = 0 
assign u[4'b1000] [59] = 22'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = 0 
assign u[4'b1000] [60] = 22'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = 0 
assign u[4'b1000] [61] = 22'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = 0 
assign u[4'b1000] [62] = 22'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = 0 
assign u[4'b1000] [63] = 22'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = 0 
assign u[4'b1000] [64] = 22'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = 0 
assign u[4'b1001] [01] = 22'h 00019F;  // +1.6218604324326575 = 2^ 1 * ln( 1 +  1 * 2^(- 1+1) + ( 1^2+ 0^2) * 2^(-2* 1) )   n =  1   d_n = 1 
assign u[4'b1001] [02] = 22'h 0001C8;  // +1.7851484105136781 = 2^ 2 * ln( 1 +  1 * 2^(- 2+1) + ( 1^2+ 0^2) * 2^(-2* 2) )   n =  2   d_n = 1 
assign u[4'b1001] [03] = 22'h 0001E2;  // +1.8845285705021353 = 2^ 3 * ln( 1 +  1 * 2^(- 3+1) + ( 1^2+ 0^2) * 2^(-2* 3) )   n =  3   d_n = 1 
assign u[4'b1001] [04] = 22'h 0001F0;  // +1.9399878981259149 = 2^ 4 * ln( 1 +  1 * 2^(- 4+1) + ( 1^2+ 0^2) * 2^(-2* 4) )   n =  4   d_n = 1 
assign u[4'b1001] [05] = 22'h 0001F8;  // +1.9693861546722360 = 2^ 5 * ln( 1 +  1 * 2^(- 5+1) + ( 1^2+ 0^2) * 2^(-2* 5) )   n =  5   d_n = 1 
assign u[4'b1001] [06] = 22'h 0001FC;  // +1.9845358766035526 = 2^ 6 * ln( 1 +  1 * 2^(- 6+1) + ( 1^2+ 0^2) * 2^(-2* 6) )   n =  6   d_n = 1 
assign u[4'b1001] [07] = 22'h 0001FE;  // +1.9922279531660669 = 2^ 7 * ln( 1 +  1 * 2^(- 7+1) + ( 1^2+ 0^2) * 2^(-2* 7) )   n =  7   d_n = 1 
assign u[4'b1001] [08] = 22'h 0001FF;  // +1.9961038928165493 = 2^ 8 * ln( 1 +  1 * 2^(- 8+1) + ( 1^2+ 0^2) * 2^(-2* 8) )   n =  8   d_n = 1 
assign u[4'b1001] [09] = 22'h 0001FF;  // +1.9980494144120313 = 2^ 9 * ln( 1 +  1 * 2^(- 9+1) + ( 1^2+ 0^2) * 2^(-2* 9) )   n =  9   d_n = 1 
assign u[4'b1001] [10] = 22'h 0001FF;  // +1.9990240728175799 = 2^10 * ln( 1 +  1 * 2^(-10+1) + ( 1^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = 1 
assign u[4'b1001] [11] = 22'h 0001FF;  // +1.9995118776375345 = 2^11 * ln( 1 +  1 * 2^(-11+1) + ( 1^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = 1 
assign u[4'b1001] [12] = 22'h 0001FF;  // +1.9997558991041553 = 2^12 * ln( 1 +  1 * 2^(-12+1) + ( 1^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = 1 
assign u[4'b1001] [13] = 22'h 0001FF;  // +1.9998779396206980 = 2^13 * ln( 1 +  1 * 2^(-13+1) + ( 1^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = 1 
assign u[4'b1001] [14] = 22'h 0001FF;  // +1.9999389673271633 = 2^14 * ln( 1 +  1 * 2^(-14+1) + ( 1^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = 1 
assign u[4'b1001] [15] = 22'h 0001FF;  // +1.9999694830427426 = 2^15 * ln( 1 +  1 * 2^(-15+1) + ( 1^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = 1 
assign u[4'b1001] [16] = 22'h 0001FF;  // +1.9999847413661562 = 2^16 * ln( 1 +  1 * 2^(-16+1) + ( 1^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = 1 
assign u[4'b1001] [17] = 22'h 0001FF;  // +1.9999923706442737 = 2^17 * ln( 1 +  1 * 2^(-17+1) + ( 1^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = 1 
assign u[4'b1001] [18] = 22'h 0001FF;  // +1.9999961853124357 = 2^18 * ln( 1 +  1 * 2^(-18+1) + ( 1^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = 1 
assign u[4'b1001] [19] = 22'h 0001FF;  // +1.9999980926537926 = 2^19 * ln( 1 +  1 * 2^(-19+1) + ( 1^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = 1 
assign u[4'b1001] [20] = 22'h 0001FF;  // +1.9999990463262900 = 2^20 * ln( 1 +  1 * 2^(-20+1) + ( 1^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = 1 
assign u[4'b1001] [21] = 22'h 0001FF;  // +1.9999995231629935 = 2^21 * ln( 1 +  1 * 2^(-21+1) + ( 1^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = 1 
assign u[4'b1001] [22] = 22'h 0001FF;  // +1.9999997615814589 = 2^22 * ln( 1 +  1 * 2^(-22+1) + ( 1^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = 1 
assign u[4'b1001] [23] = 22'h 0001FF;  // +1.9999998807907200 = 2^23 * ln( 1 +  1 * 2^(-23+1) + ( 1^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = 1 
assign u[4'b1001] [24] = 22'h 0001FF;  // +1.9999999403953577 = 2^24 * ln( 1 +  1 * 2^(-24+1) + ( 1^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = 1 
assign u[4'b1001] [25] = 22'h 0001FF;  // +1.9999999701976783 = 2^25 * ln( 1 +  1 * 2^(-25+1) + ( 1^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = 1 
assign u[4'b1001] [26] = 22'h 0001FF;  // +1.9999999850988390 = 2^26 * ln( 1 +  1 * 2^(-26+1) + ( 1^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = 1 
assign u[4'b1001] [27] = 22'h 0001FF;  // +1.9999999925494194 = 2^27 * ln( 1 +  1 * 2^(-27+1) + ( 1^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = 1 
assign u[4'b1001] [28] = 22'h 0001FF;  // +1.9999999962747097 = 2^28 * ln( 1 +  1 * 2^(-28+1) + ( 1^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = 1 
assign u[4'b1001] [29] = 22'h 0001FF;  // +1.9999999981373549 = 2^29 * ln( 1 +  1 * 2^(-29+1) + ( 1^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = 1 
assign u[4'b1001] [30] = 22'h 0001FF;  // +1.9999999990686774 = 2^30 * ln( 1 +  1 * 2^(-30+1) + ( 1^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = 1 
assign u[4'b1001] [31] = 22'h 0001FF;  // +1.9999999995343387 = 2^31 * ln( 1 +  1 * 2^(-31+1) + ( 1^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = 1 
assign u[4'b1001] [32] = 22'h 0001FF;  // +1.9999999997671694 = 2^32 * ln( 1 +  1 * 2^(-32+1) + ( 1^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = 1 
assign u[4'b1001] [33] = 22'h 0001FF;  // +1.9999999998835847 = 2^33 * ln( 1 +  1 * 2^(-33+1) + ( 1^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = 1 
assign u[4'b1001] [34] = 22'h 0001FF;  // +1.9999999999417923 = 2^34 * ln( 1 +  1 * 2^(-34+1) + ( 1^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = 1 
assign u[4'b1001] [35] = 22'h 0001FF;  // +1.9999999999708962 = 2^35 * ln( 1 +  1 * 2^(-35+1) + ( 1^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = 1 
assign u[4'b1001] [36] = 22'h 0001FF;  // +1.9999999999854481 = 2^36 * ln( 1 +  1 * 2^(-36+1) + ( 1^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = 1 
assign u[4'b1001] [37] = 22'h 0001FF;  // +1.9999999999927240 = 2^37 * ln( 1 +  1 * 2^(-37+1) + ( 1^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = 1 
assign u[4'b1001] [38] = 22'h 0001FF;  // +1.9999999999963620 = 2^38 * ln( 1 +  1 * 2^(-38+1) + ( 1^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = 1 
assign u[4'b1001] [39] = 22'h 0001FF;  // +1.9999999999981810 = 2^39 * ln( 1 +  1 * 2^(-39+1) + ( 1^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = 1 
assign u[4'b1001] [40] = 22'h 0001FF;  // +1.9999999999990905 = 2^40 * ln( 1 +  1 * 2^(-40+1) + ( 1^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = 1 
assign u[4'b1001] [41] = 22'h 0001FF;  // +1.9999999999995453 = 2^41 * ln( 1 +  1 * 2^(-41+1) + ( 1^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = 1 
assign u[4'b1001] [42] = 22'h 0001FF;  // +1.9999999999997726 = 2^42 * ln( 1 +  1 * 2^(-42+1) + ( 1^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = 1 
assign u[4'b1001] [43] = 22'h 0001FF;  // +1.9999999999998863 = 2^43 * ln( 1 +  1 * 2^(-43+1) + ( 1^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = 1 
assign u[4'b1001] [44] = 22'h 0001FF;  // +1.9999999999999432 = 2^44 * ln( 1 +  1 * 2^(-44+1) + ( 1^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = 1 
assign u[4'b1001] [45] = 22'h 0001FF;  // +1.9999999999999716 = 2^45 * ln( 1 +  1 * 2^(-45+1) + ( 1^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = 1 
assign u[4'b1001] [46] = 22'h 0001FF;  // +1.9999999999999858 = 2^46 * ln( 1 +  1 * 2^(-46+1) + ( 1^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = 1 
assign u[4'b1001] [47] = 22'h 0001FF;  // +1.9999999999999929 = 2^47 * ln( 1 +  1 * 2^(-47+1) + ( 1^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = 1 
assign u[4'b1001] [48] = 22'h 0001FF;  // +1.9999999999999964 = 2^48 * ln( 1 +  1 * 2^(-48+1) + ( 1^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = 1 
assign u[4'b1001] [49] = 22'h 0001FF;  // +1.9999999999999982 = 2^49 * ln( 1 +  1 * 2^(-49+1) + ( 1^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = 1 
assign u[4'b1001] [50] = 22'h 0001FF;  // +1.9999999999999991 = 2^50 * ln( 1 +  1 * 2^(-50+1) + ( 1^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = 1 
assign u[4'b1001] [51] = 22'h 0001FF;  // +1.9999999999999996 = 2^51 * ln( 1 +  1 * 2^(-51+1) + ( 1^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = 1 
assign u[4'b1001] [52] = 22'h 0001FF;  // +1.9999999999999998 = 2^52 * ln( 1 +  1 * 2^(-52+1) + ( 1^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = 1 
assign u[4'b1001] [53] = 22'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  1 * 2^(-53+1) + ( 1^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = 1 
assign u[4'b1001] [54] = 22'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  1 * 2^(-54+1) + ( 1^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = 1 
assign u[4'b1001] [55] = 22'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  1 * 2^(-55+1) + ( 1^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = 1 
assign u[4'b1001] [56] = 22'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  1 * 2^(-56+1) + ( 1^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = 1 
assign u[4'b1001] [57] = 22'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  1 * 2^(-57+1) + ( 1^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = 1 
assign u[4'b1001] [58] = 22'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  1 * 2^(-58+1) + ( 1^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = 1 
assign u[4'b1001] [59] = 22'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  1 * 2^(-59+1) + ( 1^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = 1 
assign u[4'b1001] [60] = 22'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  1 * 2^(-60+1) + ( 1^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = 1 
assign u[4'b1001] [61] = 22'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  1 * 2^(-61+1) + ( 1^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = 1 
assign u[4'b1001] [62] = 22'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  1 * 2^(-62+1) + ( 1^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = 1 
assign u[4'b1001] [63] = 22'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  1 * 2^(-63+1) + ( 1^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = 1 
assign u[4'b1001] [64] = 22'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  1 * 2^(-64+1) + ( 1^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = 1 
assign u[4'b1010] [01] = 22'h 000000;  // +0.0000000000000000 = 2^ 1 * ln( 1 +  0 * 2^(- 1+1) + ( 0^2+ 0^2) * 2^(-2* 1) )   n =  1   d_n = -0 
assign u[4'b1010] [02] = 22'h 000000;  // +0.0000000000000000 = 2^ 2 * ln( 1 +  0 * 2^(- 2+1) + ( 0^2+ 0^2) * 2^(-2* 2) )   n =  2   d_n = -0 
assign u[4'b1010] [03] = 22'h 000000;  // +0.0000000000000000 = 2^ 3 * ln( 1 +  0 * 2^(- 3+1) + ( 0^2+ 0^2) * 2^(-2* 3) )   n =  3   d_n = -0 
assign u[4'b1010] [04] = 22'h 000000;  // +0.0000000000000000 = 2^ 4 * ln( 1 +  0 * 2^(- 4+1) + ( 0^2+ 0^2) * 2^(-2* 4) )   n =  4   d_n = -0 
assign u[4'b1010] [05] = 22'h 000000;  // +0.0000000000000000 = 2^ 5 * ln( 1 +  0 * 2^(- 5+1) + ( 0^2+ 0^2) * 2^(-2* 5) )   n =  5   d_n = -0 
assign u[4'b1010] [06] = 22'h 000000;  // +0.0000000000000000 = 2^ 6 * ln( 1 +  0 * 2^(- 6+1) + ( 0^2+ 0^2) * 2^(-2* 6) )   n =  6   d_n = -0 
assign u[4'b1010] [07] = 22'h 000000;  // +0.0000000000000000 = 2^ 7 * ln( 1 +  0 * 2^(- 7+1) + ( 0^2+ 0^2) * 2^(-2* 7) )   n =  7   d_n = -0 
assign u[4'b1010] [08] = 22'h 000000;  // +0.0000000000000000 = 2^ 8 * ln( 1 +  0 * 2^(- 8+1) + ( 0^2+ 0^2) * 2^(-2* 8) )   n =  8   d_n = -0 
assign u[4'b1010] [09] = 22'h 000000;  // +0.0000000000000000 = 2^ 9 * ln( 1 +  0 * 2^(- 9+1) + ( 0^2+ 0^2) * 2^(-2* 9) )   n =  9   d_n = -0 
assign u[4'b1010] [10] = 22'h 000000;  // +0.0000000000000000 = 2^10 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = -0 
assign u[4'b1010] [11] = 22'h 000000;  // +0.0000000000000000 = 2^11 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = -0 
assign u[4'b1010] [12] = 22'h 000000;  // +0.0000000000000000 = 2^12 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = -0 
assign u[4'b1010] [13] = 22'h 000000;  // +0.0000000000000000 = 2^13 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = -0 
assign u[4'b1010] [14] = 22'h 000000;  // +0.0000000000000000 = 2^14 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = -0 
assign u[4'b1010] [15] = 22'h 000000;  // +0.0000000000000000 = 2^15 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = -0 
assign u[4'b1010] [16] = 22'h 000000;  // +0.0000000000000000 = 2^16 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = -0 
assign u[4'b1010] [17] = 22'h 000000;  // +0.0000000000000000 = 2^17 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = -0 
assign u[4'b1010] [18] = 22'h 000000;  // +0.0000000000000000 = 2^18 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = -0 
assign u[4'b1010] [19] = 22'h 000000;  // +0.0000000000000000 = 2^19 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = -0 
assign u[4'b1010] [20] = 22'h 000000;  // +0.0000000000000000 = 2^20 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = -0 
assign u[4'b1010] [21] = 22'h 000000;  // +0.0000000000000000 = 2^21 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = -0 
assign u[4'b1010] [22] = 22'h 000000;  // +0.0000000000000000 = 2^22 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = -0 
assign u[4'b1010] [23] = 22'h 000000;  // +0.0000000000000000 = 2^23 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = -0 
assign u[4'b1010] [24] = 22'h 000000;  // +0.0000000000000000 = 2^24 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = -0 
assign u[4'b1010] [25] = 22'h 000000;  // +0.0000000000000000 = 2^25 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = -0 
assign u[4'b1010] [26] = 22'h 000000;  // +0.0000000000000000 = 2^26 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = -0 
assign u[4'b1010] [27] = 22'h 000000;  // +0.0000000000000000 = 2^27 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = -0 
assign u[4'b1010] [28] = 22'h 000000;  // +0.0000000000000000 = 2^28 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = -0 
assign u[4'b1010] [29] = 22'h 000000;  // +0.0000000000000000 = 2^29 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = -0 
assign u[4'b1010] [30] = 22'h 000000;  // +0.0000000000000000 = 2^30 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = -0 
assign u[4'b1010] [31] = 22'h 000000;  // +0.0000000000000000 = 2^31 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = -0 
assign u[4'b1010] [32] = 22'h 000000;  // +0.0000000000000000 = 2^32 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = -0 
assign u[4'b1010] [33] = 22'h 000000;  // +0.0000000000000000 = 2^33 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = -0 
assign u[4'b1010] [34] = 22'h 000000;  // +0.0000000000000000 = 2^34 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = -0 
assign u[4'b1010] [35] = 22'h 000000;  // +0.0000000000000000 = 2^35 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = -0 
assign u[4'b1010] [36] = 22'h 000000;  // +0.0000000000000000 = 2^36 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = -0 
assign u[4'b1010] [37] = 22'h 000000;  // +0.0000000000000000 = 2^37 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = -0 
assign u[4'b1010] [38] = 22'h 000000;  // +0.0000000000000000 = 2^38 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = -0 
assign u[4'b1010] [39] = 22'h 000000;  // +0.0000000000000000 = 2^39 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = -0 
assign u[4'b1010] [40] = 22'h 000000;  // +0.0000000000000000 = 2^40 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = -0 
assign u[4'b1010] [41] = 22'h 000000;  // +0.0000000000000000 = 2^41 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = -0 
assign u[4'b1010] [42] = 22'h 000000;  // +0.0000000000000000 = 2^42 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = -0 
assign u[4'b1010] [43] = 22'h 000000;  // +0.0000000000000000 = 2^43 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = -0 
assign u[4'b1010] [44] = 22'h 000000;  // +0.0000000000000000 = 2^44 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = -0 
assign u[4'b1010] [45] = 22'h 000000;  // +0.0000000000000000 = 2^45 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = -0 
assign u[4'b1010] [46] = 22'h 000000;  // +0.0000000000000000 = 2^46 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = -0 
assign u[4'b1010] [47] = 22'h 000000;  // +0.0000000000000000 = 2^47 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = -0 
assign u[4'b1010] [48] = 22'h 000000;  // +0.0000000000000000 = 2^48 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = -0 
assign u[4'b1010] [49] = 22'h 000000;  // +0.0000000000000000 = 2^49 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = -0 
assign u[4'b1010] [50] = 22'h 000000;  // +0.0000000000000000 = 2^50 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = -0 
assign u[4'b1010] [51] = 22'h 000000;  // +0.0000000000000000 = 2^51 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = -0 
assign u[4'b1010] [52] = 22'h 000000;  // +0.0000000000000000 = 2^52 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = -0 
assign u[4'b1010] [53] = 22'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = -0 
assign u[4'b1010] [54] = 22'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = -0 
assign u[4'b1010] [55] = 22'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = -0 
assign u[4'b1010] [56] = 22'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = -0 
assign u[4'b1010] [57] = 22'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = -0 
assign u[4'b1010] [58] = 22'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = -0 
assign u[4'b1010] [59] = 22'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = -0 
assign u[4'b1010] [60] = 22'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = -0 
assign u[4'b1010] [61] = 22'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = -0 
assign u[4'b1010] [62] = 22'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = -0 
assign u[4'b1010] [63] = 22'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = -0 
assign u[4'b1010] [64] = 22'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = -0 
assign u[4'b1011] [01] = 22'h 3FFD3A;  // -2.7725887222397811 = 2^ 1 * ln( 1 + -1 * 2^(- 1+1) + (-1^2+ 0^2) * 2^(-2* 1) )   n =  1   d_n = -1 
assign u[4'b1011] [02] = 22'h 3FFDB2;  // -2.3014565796142472 = 2^ 2 * ln( 1 + -1 * 2^(- 2+1) + (-1^2+ 0^2) * 2^(-2* 2) )   n =  2   d_n = -1 
assign u[4'b1011] [03] = 22'h 3FFDDD;  // -2.1365022819923620 = 2^ 3 * ln( 1 + -1 * 2^(- 3+1) + (-1^2+ 0^2) * 2^(-2* 3) )   n =  3   d_n = -1 
assign u[4'b1011] [04] = 22'h 3FFDEF;  // -2.0652326764022777 = 2^ 4 * ln( 1 + -1 * 2^(- 4+1) + (-1^2+ 0^2) * 2^(-2* 4) )   n =  4   d_n = -1 
assign u[4'b1011] [05] = 22'h 3FFDF7;  // -2.0319166921331391 = 2^ 5 * ln( 1 + -1 * 2^(- 5+1) + (-1^2+ 0^2) * 2^(-2* 5) )   n =  5   d_n = -1 
assign u[4'b1011] [06] = 22'h 3FFDFB;  // -2.0157896919218135 = 2^ 6 * ln( 1 + -1 * 2^(- 6+1) + (-1^2+ 0^2) * 2^(-2* 6) )   n =  6   d_n = -1 
assign u[4'b1011] [07] = 22'h 3FFDFD;  // -2.0078534300226285 = 2^ 7 * ln( 1 + -1 * 2^(- 7+1) + (-1^2+ 0^2) * 2^(-2* 7) )   n =  7   d_n = -1 
assign u[4'b1011] [08] = 22'h 3FFDFE;  // -2.0039164524218003 = 2^ 8 * ln( 1 + -1 * 2^(- 8+1) + (-1^2+ 0^2) * 2^(-2* 8) )   n =  8   d_n = -1 
assign u[4'b1011] [09] = 22'h 3FFDFF;  // -2.0019556718626310 = 2^ 9 * ln( 1 + -1 * 2^(- 9+1) + (-1^2+ 0^2) * 2^(-2* 9) )   n =  9   d_n = -1 
assign u[4'b1011] [10] = 22'h 3FFDFF;  // -2.0009771987489029 = 2^10 * ln( 1 + -1 * 2^(-10+1) + (-1^2+ 0^2) * 2^(-2*10) )   n = 10   d_n = -1 
assign u[4'b1011] [11] = 22'h 3FFDFF;  // -2.0004884402539500 = 2^11 * ln( 1 + -1 * 2^(-11+1) + (-1^2+ 0^2) * 2^(-2*11) )   n = 11   d_n = -1 
assign u[4'b1011] [12] = 22'h 3FFDFF;  // -2.0002441803687074 = 2^12 * ln( 1 + -1 * 2^(-12+1) + (-1^2+ 0^2) * 2^(-2*12) )   n = 12   d_n = -1 
assign u[4'b1011] [13] = 22'h 3FFDFF;  // -2.0001220802475173 = 2^13 * ln( 1 + -1 * 2^(-13+1) + (-1^2+ 0^2) * 2^(-2*13) )   n = 13   d_n = -1 
assign u[4'b1011] [14] = 22'h 3FFDFF;  // -2.0000610376398904 = 2^14 * ln( 1 + -1 * 2^(-14+1) + (-1^2+ 0^2) * 2^(-2*14) )   n = 14   d_n = -1 
assign u[4'b1011] [15] = 22'h 3FFDFF;  // -2.0000305181990208 = 2^15 * ln( 1 + -1 * 2^(-15+1) + (-1^2+ 0^2) * 2^(-2*15) )   n = 15   d_n = -1 
assign u[4'b1011] [16] = 22'h 3FFDFF;  // -2.0000152589442846 = 2^16 * ln( 1 + -1 * 2^(-16+1) + (-1^2+ 0^2) * 2^(-2*16) )   n = 16   d_n = -1 
assign u[4'b1011] [17] = 22'h 3FFDFF;  // -2.0000076294333367 = 2^17 * ln( 1 + -1 * 2^(-17+1) + (-1^2+ 0^2) * 2^(-2*17) )   n = 17   d_n = -1 
assign u[4'b1011] [18] = 22'h 3FFDFF;  // -2.0000038147069668 = 2^18 * ln( 1 + -1 * 2^(-18+1) + (-1^2+ 0^2) * 2^(-2*18) )   n = 18   d_n = -1 
assign u[4'b1011] [19] = 22'h 3FFDFF;  // -2.0000019073510580 = 2^19 * ln( 1 + -1 * 2^(-19+1) + (-1^2+ 0^2) * 2^(-2*19) )   n = 19   d_n = -1 
assign u[4'b1011] [20] = 22'h 3FFDFF;  // -2.0000009536749226 = 2^20 * ln( 1 + -1 * 2^(-20+1) + (-1^2+ 0^2) * 2^(-2*20) )   n = 20   d_n = -1 
assign u[4'b1011] [21] = 22'h 3FFDFF;  // -2.0000004768373096 = 2^21 * ln( 1 + -1 * 2^(-21+1) + (-1^2+ 0^2) * 2^(-2*21) )   n = 21   d_n = -1 
assign u[4'b1011] [22] = 22'h 3FFDFF;  // -2.0000002384186168 = 2^22 * ln( 1 + -1 * 2^(-22+1) + (-1^2+ 0^2) * 2^(-2*22) )   n = 22   d_n = -1 
assign u[4'b1011] [23] = 22'h 3FFDFF;  // -2.0000001192092989 = 2^23 * ln( 1 + -1 * 2^(-23+1) + (-1^2+ 0^2) * 2^(-2*23) )   n = 23   d_n = -1 
assign u[4'b1011] [24] = 22'h 3FFDFF;  // -2.0000000596046470 = 2^24 * ln( 1 + -1 * 2^(-24+1) + (-1^2+ 0^2) * 2^(-2*24) )   n = 24   d_n = -1 
assign u[4'b1011] [25] = 22'h 3FFDFF;  // -2.0000000298023228 = 2^25 * ln( 1 + -1 * 2^(-25+1) + (-1^2+ 0^2) * 2^(-2*25) )   n = 25   d_n = -1 
assign u[4'b1011] [26] = 22'h 3FFDFF;  // -2.0000000149011612 = 2^26 * ln( 1 + -1 * 2^(-26+1) + (-1^2+ 0^2) * 2^(-2*26) )   n = 26   d_n = -1 
assign u[4'b1011] [27] = 22'h 3FFDFF;  // -2.0000000074505806 = 2^27 * ln( 1 + -1 * 2^(-27+1) + (-1^2+ 0^2) * 2^(-2*27) )   n = 27   d_n = -1 
assign u[4'b1011] [28] = 22'h 3FFDFF;  // -2.0000000037252903 = 2^28 * ln( 1 + -1 * 2^(-28+1) + (-1^2+ 0^2) * 2^(-2*28) )   n = 28   d_n = -1 
assign u[4'b1011] [29] = 22'h 3FFDFF;  // -2.0000000018626451 = 2^29 * ln( 1 + -1 * 2^(-29+1) + (-1^2+ 0^2) * 2^(-2*29) )   n = 29   d_n = -1 
assign u[4'b1011] [30] = 22'h 3FFDFF;  // -2.0000000009313226 = 2^30 * ln( 1 + -1 * 2^(-30+1) + (-1^2+ 0^2) * 2^(-2*30) )   n = 30   d_n = -1 
assign u[4'b1011] [31] = 22'h 3FFDFF;  // -2.0000000004656613 = 2^31 * ln( 1 + -1 * 2^(-31+1) + (-1^2+ 0^2) * 2^(-2*31) )   n = 31   d_n = -1 
assign u[4'b1011] [32] = 22'h 3FFDFF;  // -2.0000000002328306 = 2^32 * ln( 1 + -1 * 2^(-32+1) + (-1^2+ 0^2) * 2^(-2*32) )   n = 32   d_n = -1 
assign u[4'b1011] [33] = 22'h 3FFDFF;  // -2.0000000001164153 = 2^33 * ln( 1 + -1 * 2^(-33+1) + (-1^2+ 0^2) * 2^(-2*33) )   n = 33   d_n = -1 
assign u[4'b1011] [34] = 22'h 3FFDFF;  // -2.0000000000582077 = 2^34 * ln( 1 + -1 * 2^(-34+1) + (-1^2+ 0^2) * 2^(-2*34) )   n = 34   d_n = -1 
assign u[4'b1011] [35] = 22'h 3FFDFF;  // -2.0000000000291038 = 2^35 * ln( 1 + -1 * 2^(-35+1) + (-1^2+ 0^2) * 2^(-2*35) )   n = 35   d_n = -1 
assign u[4'b1011] [36] = 22'h 3FFDFF;  // -2.0000000000145519 = 2^36 * ln( 1 + -1 * 2^(-36+1) + (-1^2+ 0^2) * 2^(-2*36) )   n = 36   d_n = -1 
assign u[4'b1011] [37] = 22'h 3FFDFF;  // -2.0000000000072760 = 2^37 * ln( 1 + -1 * 2^(-37+1) + (-1^2+ 0^2) * 2^(-2*37) )   n = 37   d_n = -1 
assign u[4'b1011] [38] = 22'h 3FFDFF;  // -2.0000000000036380 = 2^38 * ln( 1 + -1 * 2^(-38+1) + (-1^2+ 0^2) * 2^(-2*38) )   n = 38   d_n = -1 
assign u[4'b1011] [39] = 22'h 3FFDFF;  // -2.0000000000018190 = 2^39 * ln( 1 + -1 * 2^(-39+1) + (-1^2+ 0^2) * 2^(-2*39) )   n = 39   d_n = -1 
assign u[4'b1011] [40] = 22'h 3FFE00;  // -2.0000000000009095 = 2^40 * ln( 1 + -1 * 2^(-40+1) + (-1^2+ 0^2) * 2^(-2*40) )   n = 40   d_n = -1 
assign u[4'b1011] [41] = 22'h 3FFE00;  // -2.0000000000004547 = 2^41 * ln( 1 + -1 * 2^(-41+1) + (-1^2+ 0^2) * 2^(-2*41) )   n = 41   d_n = -1 
assign u[4'b1011] [42] = 22'h 3FFE00;  // -2.0000000000002274 = 2^42 * ln( 1 + -1 * 2^(-42+1) + (-1^2+ 0^2) * 2^(-2*42) )   n = 42   d_n = -1 
assign u[4'b1011] [43] = 22'h 3FFE00;  // -2.0000000000001137 = 2^43 * ln( 1 + -1 * 2^(-43+1) + (-1^2+ 0^2) * 2^(-2*43) )   n = 43   d_n = -1 
assign u[4'b1011] [44] = 22'h 3FFE00;  // -2.0000000000000568 = 2^44 * ln( 1 + -1 * 2^(-44+1) + (-1^2+ 0^2) * 2^(-2*44) )   n = 44   d_n = -1 
assign u[4'b1011] [45] = 22'h 3FFE00;  // -2.0000000000000284 = 2^45 * ln( 1 + -1 * 2^(-45+1) + (-1^2+ 0^2) * 2^(-2*45) )   n = 45   d_n = -1 
assign u[4'b1011] [46] = 22'h 3FFE00;  // -2.0000000000000142 = 2^46 * ln( 1 + -1 * 2^(-46+1) + (-1^2+ 0^2) * 2^(-2*46) )   n = 46   d_n = -1 
assign u[4'b1011] [47] = 22'h 3FFE00;  // -2.0000000000000071 = 2^47 * ln( 1 + -1 * 2^(-47+1) + (-1^2+ 0^2) * 2^(-2*47) )   n = 47   d_n = -1 
assign u[4'b1011] [48] = 22'h 3FFE00;  // -2.0000000000000036 = 2^48 * ln( 1 + -1 * 2^(-48+1) + (-1^2+ 0^2) * 2^(-2*48) )   n = 48   d_n = -1 
assign u[4'b1011] [49] = 22'h 3FFE00;  // -2.0000000000000018 = 2^49 * ln( 1 + -1 * 2^(-49+1) + (-1^2+ 0^2) * 2^(-2*49) )   n = 49   d_n = -1 
assign u[4'b1011] [50] = 22'h 3FFE00;  // -2.0000000000000009 = 2^50 * ln( 1 + -1 * 2^(-50+1) + (-1^2+ 0^2) * 2^(-2*50) )   n = 50   d_n = -1 
assign u[4'b1011] [51] = 22'h 3FFE00;  // -2.0000000000000004 = 2^51 * ln( 1 + -1 * 2^(-51+1) + (-1^2+ 0^2) * 2^(-2*51) )   n = 51   d_n = -1 
assign u[4'b1011] [52] = 22'h 3FFE00;  // -2.0000000000000004 = 2^52 * ln( 1 + -1 * 2^(-52+1) + (-1^2+ 0^2) * 2^(-2*52) )   n = 52   d_n = -1 
assign u[4'b1011] [53] = 22'h 3FFE00;  // -2.0000000000000000 = 2^53 * ln( 1 + -1 * 2^(-53+1) + (-1^2+ 0^2) * 2^(-2*53) )   n = 53   d_n = -1 
assign u[4'b1011] [54] = 22'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 + -1 * 2^(-54+1) + (-1^2+ 0^2) * 2^(-2*54) )   n = 54   d_n = -1 
assign u[4'b1011] [55] = 22'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 + -1 * 2^(-55+1) + (-1^2+ 0^2) * 2^(-2*55) )   n = 55   d_n = -1 
assign u[4'b1011] [56] = 22'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 + -1 * 2^(-56+1) + (-1^2+ 0^2) * 2^(-2*56) )   n = 56   d_n = -1 
assign u[4'b1011] [57] = 22'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 + -1 * 2^(-57+1) + (-1^2+ 0^2) * 2^(-2*57) )   n = 57   d_n = -1 
assign u[4'b1011] [58] = 22'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 + -1 * 2^(-58+1) + (-1^2+ 0^2) * 2^(-2*58) )   n = 58   d_n = -1 
assign u[4'b1011] [59] = 22'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 + -1 * 2^(-59+1) + (-1^2+ 0^2) * 2^(-2*59) )   n = 59   d_n = -1 
assign u[4'b1011] [60] = 22'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 + -1 * 2^(-60+1) + (-1^2+ 0^2) * 2^(-2*60) )   n = 60   d_n = -1 
assign u[4'b1011] [61] = 22'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 + -1 * 2^(-61+1) + (-1^2+ 0^2) * 2^(-2*61) )   n = 61   d_n = -1 
assign u[4'b1011] [62] = 22'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 + -1 * 2^(-62+1) + (-1^2+ 0^2) * 2^(-2*62) )   n = 62   d_n = -1 
assign u[4'b1011] [63] = 22'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 + -1 * 2^(-63+1) + (-1^2+ 0^2) * 2^(-2*63) )   n = 63   d_n = -1 
assign u[4'b1011] [64] = 22'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 + -1 * 2^(-64+1) + (-1^2+ 0^2) * 2^(-2*64) )   n = 64   d_n = -1 
assign u[4'b1100] [01] = 22'h 000072;  // +0.4462871026284197 = 2^ 1 * ln( 1 +  0 * 2^(- 1+1) + ( 0^2+-1^2) * 2^(-2* 1) )   n =  1   d_n = -0-1i 
assign u[4'b1100] [02] = 22'h 00003E;  // +0.2424984872657394 = 2^ 2 * ln( 1 +  0 * 2^(- 2+1) + ( 0^2+-1^2) * 2^(-2* 2) )   n =  2   d_n = -0-1i 
assign u[4'b1100] [03] = 22'h 00001F;  // +0.1240334922877210 = 2^ 3 * ln( 1 +  0 * 2^(- 3+1) + ( 0^2+-1^2) * 2^(-2* 3) )   n =  3   d_n = -0-1i 
assign u[4'b1100] [04] = 22'h 00000F;  // +0.0623782466505195 = 2^ 4 * ln( 1 +  0 * 2^(- 4+1) + ( 0^2+-1^2) * 2^(-2* 4) )   n =  4   d_n = -0-1i 
assign u[4'b1100] [05] = 22'h 000007;  // +0.0312347511377731 = 2^ 5 * ln( 1 +  0 * 2^(- 5+1) + ( 0^2+-1^2) * 2^(-2* 5) )   n =  5   d_n = -0-1i 
assign u[4'b1100] [06] = 22'h 000003;  // +0.0156230929617406 = 2^ 6 * ln( 1 +  0 * 2^(- 6+1) + ( 0^2+-1^2) * 2^(-2* 6) )   n =  6   d_n = -0-1i 
assign u[4'b1100] [07] = 22'h 000001;  // +0.0078122615911219 = 2^ 7 * ln( 1 +  0 * 2^(- 7+1) + ( 0^2+-1^2) * 2^(-2* 7) )   n =  7   d_n = -0-1i 
assign u[4'b1100] [08] = 22'h 000000;  // +0.0039062201979808 = 2^ 8 * ln( 1 +  0 * 2^(- 8+1) + ( 0^2+-1^2) * 2^(-2* 8) )   n =  8   d_n = -0-1i 
assign u[4'b1100] [09] = 22'h 000000;  // +0.0019531212747156 = 2^ 9 * ln( 1 +  0 * 2^(- 9+1) + ( 0^2+-1^2) * 2^(-2* 9) )   n =  9   d_n = -0-1i 
assign u[4'b1100] [10] = 22'h 000000;  // +0.0009765620343389 = 2^10 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+-1^2) * 2^(-2*10) )   n = 10   d_n = -0-1i 
assign u[4'b1100] [11] = 22'h 000000;  // +0.0004882811917923 = 2^11 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+-1^2) * 2^(-2*11) )   n = 11   d_n = -0-1i 
assign u[4'b1100] [12] = 22'h 000000;  // +0.0002441406177240 = 2^12 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+-1^2) * 2^(-2*12) )   n = 12   d_n = -0-1i 
assign u[4'b1100] [13] = 22'h 000000;  // +0.0001220703120453 = 2^13 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+-1^2) * 2^(-2*13) )   n = 13   d_n = -0-1i 
assign u[4'b1100] [14] = 22'h 000000;  // +0.0000610351561932 = 2^14 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+-1^2) * 2^(-2*14) )   n = 14   d_n = -0-1i 
assign u[4'b1100] [15] = 22'h 000000;  // +0.0000305175781179 = 2^15 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+-1^2) * 2^(-2*15) )   n = 15   d_n = -0-1i 
assign u[4'b1100] [16] = 22'h 000000;  // +0.0000152587890616 = 2^16 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+-1^2) * 2^(-2*16) )   n = 16   d_n = -0-1i 
assign u[4'b1100] [17] = 22'h 000000;  // +0.0000076293945311 = 2^17 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+-1^2) * 2^(-2*17) )   n = 17   d_n = -0-1i 
assign u[4'b1100] [18] = 22'h 000000;  // +0.0000038146972656 = 2^18 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+-1^2) * 2^(-2*18) )   n = 18   d_n = -0-1i 
assign u[4'b1100] [19] = 22'h 000000;  // +0.0000019073486328 = 2^19 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+-1^2) * 2^(-2*19) )   n = 19   d_n = -0-1i 
assign u[4'b1100] [20] = 22'h 000000;  // +0.0000009536743164 = 2^20 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+-1^2) * 2^(-2*20) )   n = 20   d_n = -0-1i 
assign u[4'b1100] [21] = 22'h 000000;  // +0.0000004768371582 = 2^21 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+-1^2) * 2^(-2*21) )   n = 21   d_n = -0-1i 
assign u[4'b1100] [22] = 22'h 000000;  // +0.0000002384185791 = 2^22 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+-1^2) * 2^(-2*22) )   n = 22   d_n = -0-1i 
assign u[4'b1100] [23] = 22'h 000000;  // +0.0000001192092896 = 2^23 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+-1^2) * 2^(-2*23) )   n = 23   d_n = -0-1i 
assign u[4'b1100] [24] = 22'h 000000;  // +0.0000000596046448 = 2^24 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+-1^2) * 2^(-2*24) )   n = 24   d_n = -0-1i 
assign u[4'b1100] [25] = 22'h 000000;  // +0.0000000298023224 = 2^25 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+-1^2) * 2^(-2*25) )   n = 25   d_n = -0-1i 
assign u[4'b1100] [26] = 22'h 000000;  // +0.0000000000000000 = 2^26 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+-1^2) * 2^(-2*26) )   n = 26   d_n = -0-1i 
assign u[4'b1100] [27] = 22'h 000000;  // +0.0000000000000000 = 2^27 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+-1^2) * 2^(-2*27) )   n = 27   d_n = -0-1i 
assign u[4'b1100] [28] = 22'h 000000;  // +0.0000000000000000 = 2^28 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+-1^2) * 2^(-2*28) )   n = 28   d_n = -0-1i 
assign u[4'b1100] [29] = 22'h 000000;  // +0.0000000000000000 = 2^29 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+-1^2) * 2^(-2*29) )   n = 29   d_n = -0-1i 
assign u[4'b1100] [30] = 22'h 000000;  // +0.0000000000000000 = 2^30 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+-1^2) * 2^(-2*30) )   n = 30   d_n = -0-1i 
assign u[4'b1100] [31] = 22'h 000000;  // +0.0000000000000000 = 2^31 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+-1^2) * 2^(-2*31) )   n = 31   d_n = -0-1i 
assign u[4'b1100] [32] = 22'h 000000;  // +0.0000000000000000 = 2^32 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+-1^2) * 2^(-2*32) )   n = 32   d_n = -0-1i 
assign u[4'b1100] [33] = 22'h 000000;  // +0.0000000000000000 = 2^33 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+-1^2) * 2^(-2*33) )   n = 33   d_n = -0-1i 
assign u[4'b1100] [34] = 22'h 000000;  // +0.0000000000000000 = 2^34 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+-1^2) * 2^(-2*34) )   n = 34   d_n = -0-1i 
assign u[4'b1100] [35] = 22'h 000000;  // +0.0000000000000000 = 2^35 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+-1^2) * 2^(-2*35) )   n = 35   d_n = -0-1i 
assign u[4'b1100] [36] = 22'h 000000;  // +0.0000000000000000 = 2^36 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+-1^2) * 2^(-2*36) )   n = 36   d_n = -0-1i 
assign u[4'b1100] [37] = 22'h 000000;  // +0.0000000000000000 = 2^37 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+-1^2) * 2^(-2*37) )   n = 37   d_n = -0-1i 
assign u[4'b1100] [38] = 22'h 000000;  // +0.0000000000000000 = 2^38 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+-1^2) * 2^(-2*38) )   n = 38   d_n = -0-1i 
assign u[4'b1100] [39] = 22'h 000000;  // +0.0000000000000000 = 2^39 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+-1^2) * 2^(-2*39) )   n = 39   d_n = -0-1i 
assign u[4'b1100] [40] = 22'h 000000;  // +0.0000000000000000 = 2^40 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+-1^2) * 2^(-2*40) )   n = 40   d_n = -0-1i 
assign u[4'b1100] [41] = 22'h 000000;  // +0.0000000000000000 = 2^41 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+-1^2) * 2^(-2*41) )   n = 41   d_n = -0-1i 
assign u[4'b1100] [42] = 22'h 000000;  // +0.0000000000000000 = 2^42 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+-1^2) * 2^(-2*42) )   n = 42   d_n = -0-1i 
assign u[4'b1100] [43] = 22'h 000000;  // +0.0000000000000000 = 2^43 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+-1^2) * 2^(-2*43) )   n = 43   d_n = -0-1i 
assign u[4'b1100] [44] = 22'h 000000;  // +0.0000000000000000 = 2^44 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+-1^2) * 2^(-2*44) )   n = 44   d_n = -0-1i 
assign u[4'b1100] [45] = 22'h 000000;  // +0.0000000000000000 = 2^45 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+-1^2) * 2^(-2*45) )   n = 45   d_n = -0-1i 
assign u[4'b1100] [46] = 22'h 000000;  // +0.0000000000000000 = 2^46 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+-1^2) * 2^(-2*46) )   n = 46   d_n = -0-1i 
assign u[4'b1100] [47] = 22'h 000000;  // +0.0000000000000000 = 2^47 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+-1^2) * 2^(-2*47) )   n = 47   d_n = -0-1i 
assign u[4'b1100] [48] = 22'h 000000;  // +0.0000000000000000 = 2^48 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+-1^2) * 2^(-2*48) )   n = 48   d_n = -0-1i 
assign u[4'b1100] [49] = 22'h 000000;  // +0.0000000000000000 = 2^49 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+-1^2) * 2^(-2*49) )   n = 49   d_n = -0-1i 
assign u[4'b1100] [50] = 22'h 000000;  // +0.0000000000000000 = 2^50 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+-1^2) * 2^(-2*50) )   n = 50   d_n = -0-1i 
assign u[4'b1100] [51] = 22'h 000000;  // +0.0000000000000000 = 2^51 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+-1^2) * 2^(-2*51) )   n = 51   d_n = -0-1i 
assign u[4'b1100] [52] = 22'h 000000;  // +0.0000000000000000 = 2^52 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+-1^2) * 2^(-2*52) )   n = 52   d_n = -0-1i 
assign u[4'b1100] [53] = 22'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+-1^2) * 2^(-2*53) )   n = 53   d_n = -0-1i 
assign u[4'b1100] [54] = 22'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+-1^2) * 2^(-2*54) )   n = 54   d_n = -0-1i 
assign u[4'b1100] [55] = 22'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+-1^2) * 2^(-2*55) )   n = 55   d_n = -0-1i 
assign u[4'b1100] [56] = 22'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+-1^2) * 2^(-2*56) )   n = 56   d_n = -0-1i 
assign u[4'b1100] [57] = 22'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+-1^2) * 2^(-2*57) )   n = 57   d_n = -0-1i 
assign u[4'b1100] [58] = 22'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+-1^2) * 2^(-2*58) )   n = 58   d_n = -0-1i 
assign u[4'b1100] [59] = 22'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+-1^2) * 2^(-2*59) )   n = 59   d_n = -0-1i 
assign u[4'b1100] [60] = 22'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+-1^2) * 2^(-2*60) )   n = 60   d_n = -0-1i 
assign u[4'b1100] [61] = 22'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+-1^2) * 2^(-2*61) )   n = 61   d_n = -0-1i 
assign u[4'b1100] [62] = 22'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+-1^2) * 2^(-2*62) )   n = 62   d_n = -0-1i 
assign u[4'b1100] [63] = 22'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+-1^2) * 2^(-2*63) )   n = 63   d_n = -0-1i 
assign u[4'b1100] [64] = 22'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+-1^2) * 2^(-2*64) )   n = 64   d_n = -0-1i 
assign u[4'b1101] [01] = 22'h 0001D5;  // +1.8325814637483104 = 2^ 1 * ln( 1 +  1 * 2^(- 1+1) + ( 1^2+-1^2) * 2^(-2* 1) )   n =  1   d_n = 1-1i 
assign u[4'b1101] [02] = 22'h 0001F1;  // +1.9420312631268026 = 2^ 2 * ln( 1 +  1 * 2^(- 2+1) + ( 1^2+-1^2) * 2^(-2* 2) )   n =  2   d_n = 1-1i 
assign u[4'b1101] [03] = 22'h 0001FB;  // +1.9826893112366513 = 2^ 3 * ln( 1 +  1 * 2^(- 3+1) + ( 1^2+-1^2) * 2^(-2* 3) )   n =  3   d_n = 1-1i 
assign u[4'b1101] [04] = 22'h 0001FE;  // +1.9952556560153185 = 2^ 4 * ln( 1 +  1 * 2^(- 4+1) + ( 1^2+-1^2) * 2^(-2* 4) )   n =  4   d_n = 1-1i 
assign u[4'b1101] [05] = 22'h 0001FF;  // +1.9987574279595595 = 2^ 5 * ln( 1 +  1 * 2^(- 5+1) + ( 1^2+-1^2) * 2^(-2* 5) )   n =  5   d_n = 1-1i 
assign u[4'b1101] [06] = 22'h 0001FF;  // +1.9996820132261188 = 2^ 6 * ln( 1 +  1 * 2^(- 6+1) + ( 1^2+-1^2) * 2^(-2* 6) )   n =  6   d_n = 1-1i 
assign u[4'b1101] [07] = 22'h 0001FF;  // +1.9999195675060046 = 2^ 7 * ln( 1 +  1 * 2^(- 7+1) + ( 1^2+-1^2) * 2^(-2* 7) )   n =  7   d_n = 1-1i 
assign u[4'b1101] [08] = 22'h 0001FF;  // +1.9999797737846823 = 2^ 8 * ln( 1 +  1 * 2^(- 8+1) + ( 1^2+-1^2) * 2^(-2* 8) )   n =  8   d_n = 1-1i 
assign u[4'b1101] [09] = 22'h 0001FF;  // +1.9999949286148679 = 2^ 9 * ln( 1 +  1 * 2^(- 9+1) + ( 1^2+-1^2) * 2^(-2* 9) )   n =  9   d_n = 1-1i 
assign u[4'b1101] [10] = 22'h 0001FF;  // +1.9999987302952080 = 2^10 * ln( 1 +  1 * 2^(-10+1) + ( 1^2+-1^2) * 2^(-2*10) )   n = 10   d_n = 1-1i 
assign u[4'b1101] [11] = 22'h 0001FF;  // +1.9999996823413151 = 2^11 * ln( 1 +  1 * 2^(-11+1) + ( 1^2+-1^2) * 2^(-2*11) )   n = 11   d_n = 1-1i 
assign u[4'b1101] [12] = 22'h 0001FF;  // +1.9999999205562393 = 2^12 * ln( 1 +  1 * 2^(-12+1) + ( 1^2+-1^2) * 2^(-2*12) )   n = 12   d_n = 1-1i 
assign u[4'b1101] [13] = 22'h 0001FF;  // +1.9999999801340587 = 2^13 * ln( 1 +  1 * 2^(-13+1) + ( 1^2+-1^2) * 2^(-2*13) )   n = 13   d_n = 1-1i 
assign u[4'b1101] [14] = 22'h 0001FF;  // +1.9999999950332306 = 2^14 * ln( 1 +  1 * 2^(-14+1) + ( 1^2+-1^2) * 2^(-2*14) )   n = 14   d_n = 1-1i 
assign u[4'b1101] [15] = 22'h 0001FF;  // +1.9999999987582722 = 2^15 * ln( 1 +  1 * 2^(-15+1) + ( 1^2+-1^2) * 2^(-2*15) )   n = 15   d_n = 1-1i 
assign u[4'b1101] [16] = 22'h 0001FF;  // +1.9999999996895637 = 2^16 * ln( 1 +  1 * 2^(-16+1) + ( 1^2+-1^2) * 2^(-2*16) )   n = 16   d_n = 1-1i 
assign u[4'b1101] [17] = 22'h 0001FF;  // +1.9999999999223903 = 2^17 * ln( 1 +  1 * 2^(-17+1) + ( 1^2+-1^2) * 2^(-2*17) )   n = 17   d_n = 1-1i 
assign u[4'b1101] [18] = 22'h 0001FF;  // +1.9999999999951494 = 2^18 * ln( 1 +  1 * 2^(-18+1) + ( 1^2+-1^2) * 2^(-2*18) )   n = 18   d_n = 1-1i 
assign u[4'b1101] [19] = 22'h 0001FF;  // +1.9999999999987874 = 2^19 * ln( 1 +  1 * 2^(-19+1) + ( 1^2+-1^2) * 2^(-2*19) )   n = 19   d_n = 1-1i 
assign u[4'b1101] [20] = 22'h 0001FF;  // +1.9999999999996969 = 2^20 * ln( 1 +  1 * 2^(-20+1) + ( 1^2+-1^2) * 2^(-2*20) )   n = 20   d_n = 1-1i 
assign u[4'b1101] [21] = 22'h 0001FF;  // +1.9999999999999243 = 2^21 * ln( 1 +  1 * 2^(-21+1) + ( 1^2+-1^2) * 2^(-2*21) )   n = 21   d_n = 1-1i 
assign u[4'b1101] [22] = 22'h 0001FF;  // +1.9999999999999811 = 2^22 * ln( 1 +  1 * 2^(-22+1) + ( 1^2+-1^2) * 2^(-2*22) )   n = 22   d_n = 1-1i 
assign u[4'b1101] [23] = 22'h 0001FF;  // +1.9999999999999953 = 2^23 * ln( 1 +  1 * 2^(-23+1) + ( 1^2+-1^2) * 2^(-2*23) )   n = 23   d_n = 1-1i 
assign u[4'b1101] [24] = 22'h 0001FF;  // +1.9999999999999989 = 2^24 * ln( 1 +  1 * 2^(-24+1) + ( 1^2+-1^2) * 2^(-2*24) )   n = 24   d_n = 1-1i 
assign u[4'b1101] [25] = 22'h 0001FF;  // +1.9999999999999998 = 2^25 * ln( 1 +  1 * 2^(-25+1) + ( 1^2+-1^2) * 2^(-2*25) )   n = 25   d_n = 1-1i 
assign u[4'b1101] [26] = 22'h 0001FF;  // +1.9999999850988390 = 2^26 * ln( 1 +  1 * 2^(-26+1) + ( 1^2+-1^2) * 2^(-2*26) )   n = 26   d_n = 1-1i 
assign u[4'b1101] [27] = 22'h 0001FF;  // +1.9999999925494194 = 2^27 * ln( 1 +  1 * 2^(-27+1) + ( 1^2+-1^2) * 2^(-2*27) )   n = 27   d_n = 1-1i 
assign u[4'b1101] [28] = 22'h 0001FF;  // +1.9999999962747097 = 2^28 * ln( 1 +  1 * 2^(-28+1) + ( 1^2+-1^2) * 2^(-2*28) )   n = 28   d_n = 1-1i 
assign u[4'b1101] [29] = 22'h 0001FF;  // +1.9999999981373549 = 2^29 * ln( 1 +  1 * 2^(-29+1) + ( 1^2+-1^2) * 2^(-2*29) )   n = 29   d_n = 1-1i 
assign u[4'b1101] [30] = 22'h 0001FF;  // +1.9999999990686774 = 2^30 * ln( 1 +  1 * 2^(-30+1) + ( 1^2+-1^2) * 2^(-2*30) )   n = 30   d_n = 1-1i 
assign u[4'b1101] [31] = 22'h 0001FF;  // +1.9999999995343387 = 2^31 * ln( 1 +  1 * 2^(-31+1) + ( 1^2+-1^2) * 2^(-2*31) )   n = 31   d_n = 1-1i 
assign u[4'b1101] [32] = 22'h 0001FF;  // +1.9999999997671694 = 2^32 * ln( 1 +  1 * 2^(-32+1) + ( 1^2+-1^2) * 2^(-2*32) )   n = 32   d_n = 1-1i 
assign u[4'b1101] [33] = 22'h 0001FF;  // +1.9999999998835847 = 2^33 * ln( 1 +  1 * 2^(-33+1) + ( 1^2+-1^2) * 2^(-2*33) )   n = 33   d_n = 1-1i 
assign u[4'b1101] [34] = 22'h 0001FF;  // +1.9999999999417923 = 2^34 * ln( 1 +  1 * 2^(-34+1) + ( 1^2+-1^2) * 2^(-2*34) )   n = 34   d_n = 1-1i 
assign u[4'b1101] [35] = 22'h 0001FF;  // +1.9999999999708962 = 2^35 * ln( 1 +  1 * 2^(-35+1) + ( 1^2+-1^2) * 2^(-2*35) )   n = 35   d_n = 1-1i 
assign u[4'b1101] [36] = 22'h 0001FF;  // +1.9999999999854481 = 2^36 * ln( 1 +  1 * 2^(-36+1) + ( 1^2+-1^2) * 2^(-2*36) )   n = 36   d_n = 1-1i 
assign u[4'b1101] [37] = 22'h 0001FF;  // +1.9999999999927240 = 2^37 * ln( 1 +  1 * 2^(-37+1) + ( 1^2+-1^2) * 2^(-2*37) )   n = 37   d_n = 1-1i 
assign u[4'b1101] [38] = 22'h 0001FF;  // +1.9999999999963620 = 2^38 * ln( 1 +  1 * 2^(-38+1) + ( 1^2+-1^2) * 2^(-2*38) )   n = 38   d_n = 1-1i 
assign u[4'b1101] [39] = 22'h 0001FF;  // +1.9999999999981810 = 2^39 * ln( 1 +  1 * 2^(-39+1) + ( 1^2+-1^2) * 2^(-2*39) )   n = 39   d_n = 1-1i 
assign u[4'b1101] [40] = 22'h 0001FF;  // +1.9999999999990905 = 2^40 * ln( 1 +  1 * 2^(-40+1) + ( 1^2+-1^2) * 2^(-2*40) )   n = 40   d_n = 1-1i 
assign u[4'b1101] [41] = 22'h 0001FF;  // +1.9999999999995453 = 2^41 * ln( 1 +  1 * 2^(-41+1) + ( 1^2+-1^2) * 2^(-2*41) )   n = 41   d_n = 1-1i 
assign u[4'b1101] [42] = 22'h 0001FF;  // +1.9999999999997726 = 2^42 * ln( 1 +  1 * 2^(-42+1) + ( 1^2+-1^2) * 2^(-2*42) )   n = 42   d_n = 1-1i 
assign u[4'b1101] [43] = 22'h 0001FF;  // +1.9999999999998863 = 2^43 * ln( 1 +  1 * 2^(-43+1) + ( 1^2+-1^2) * 2^(-2*43) )   n = 43   d_n = 1-1i 
assign u[4'b1101] [44] = 22'h 0001FF;  // +1.9999999999999432 = 2^44 * ln( 1 +  1 * 2^(-44+1) + ( 1^2+-1^2) * 2^(-2*44) )   n = 44   d_n = 1-1i 
assign u[4'b1101] [45] = 22'h 0001FF;  // +1.9999999999999716 = 2^45 * ln( 1 +  1 * 2^(-45+1) + ( 1^2+-1^2) * 2^(-2*45) )   n = 45   d_n = 1-1i 
assign u[4'b1101] [46] = 22'h 0001FF;  // +1.9999999999999858 = 2^46 * ln( 1 +  1 * 2^(-46+1) + ( 1^2+-1^2) * 2^(-2*46) )   n = 46   d_n = 1-1i 
assign u[4'b1101] [47] = 22'h 0001FF;  // +1.9999999999999929 = 2^47 * ln( 1 +  1 * 2^(-47+1) + ( 1^2+-1^2) * 2^(-2*47) )   n = 47   d_n = 1-1i 
assign u[4'b1101] [48] = 22'h 0001FF;  // +1.9999999999999964 = 2^48 * ln( 1 +  1 * 2^(-48+1) + ( 1^2+-1^2) * 2^(-2*48) )   n = 48   d_n = 1-1i 
assign u[4'b1101] [49] = 22'h 0001FF;  // +1.9999999999999982 = 2^49 * ln( 1 +  1 * 2^(-49+1) + ( 1^2+-1^2) * 2^(-2*49) )   n = 49   d_n = 1-1i 
assign u[4'b1101] [50] = 22'h 0001FF;  // +1.9999999999999991 = 2^50 * ln( 1 +  1 * 2^(-50+1) + ( 1^2+-1^2) * 2^(-2*50) )   n = 50   d_n = 1-1i 
assign u[4'b1101] [51] = 22'h 0001FF;  // +1.9999999999999996 = 2^51 * ln( 1 +  1 * 2^(-51+1) + ( 1^2+-1^2) * 2^(-2*51) )   n = 51   d_n = 1-1i 
assign u[4'b1101] [52] = 22'h 0001FF;  // +1.9999999999999998 = 2^52 * ln( 1 +  1 * 2^(-52+1) + ( 1^2+-1^2) * 2^(-2*52) )   n = 52   d_n = 1-1i 
assign u[4'b1101] [53] = 22'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  1 * 2^(-53+1) + ( 1^2+-1^2) * 2^(-2*53) )   n = 53   d_n = 1-1i 
assign u[4'b1101] [54] = 22'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  1 * 2^(-54+1) + ( 1^2+-1^2) * 2^(-2*54) )   n = 54   d_n = 1-1i 
assign u[4'b1101] [55] = 22'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  1 * 2^(-55+1) + ( 1^2+-1^2) * 2^(-2*55) )   n = 55   d_n = 1-1i 
assign u[4'b1101] [56] = 22'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  1 * 2^(-56+1) + ( 1^2+-1^2) * 2^(-2*56) )   n = 56   d_n = 1-1i 
assign u[4'b1101] [57] = 22'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  1 * 2^(-57+1) + ( 1^2+-1^2) * 2^(-2*57) )   n = 57   d_n = 1-1i 
assign u[4'b1101] [58] = 22'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  1 * 2^(-58+1) + ( 1^2+-1^2) * 2^(-2*58) )   n = 58   d_n = 1-1i 
assign u[4'b1101] [59] = 22'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  1 * 2^(-59+1) + ( 1^2+-1^2) * 2^(-2*59) )   n = 59   d_n = 1-1i 
assign u[4'b1101] [60] = 22'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  1 * 2^(-60+1) + ( 1^2+-1^2) * 2^(-2*60) )   n = 60   d_n = 1-1i 
assign u[4'b1101] [61] = 22'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  1 * 2^(-61+1) + ( 1^2+-1^2) * 2^(-2*61) )   n = 61   d_n = 1-1i 
assign u[4'b1101] [62] = 22'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  1 * 2^(-62+1) + ( 1^2+-1^2) * 2^(-2*62) )   n = 62   d_n = 1-1i 
assign u[4'b1101] [63] = 22'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  1 * 2^(-63+1) + ( 1^2+-1^2) * 2^(-2*63) )   n = 63   d_n = 1-1i 
assign u[4'b1101] [64] = 22'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  1 * 2^(-64+1) + ( 1^2+-1^2) * 2^(-2*64) )   n = 64   d_n = 1-1i 
assign u[4'b1110] [01] = 22'h 000072;  // +0.4462871026284197 = 2^ 1 * ln( 1 +  0 * 2^(- 1+1) + ( 0^2+-1^2) * 2^(-2* 1) )   n =  1   d_n = -0-1i 
assign u[4'b1110] [02] = 22'h 00003E;  // +0.2424984872657394 = 2^ 2 * ln( 1 +  0 * 2^(- 2+1) + ( 0^2+-1^2) * 2^(-2* 2) )   n =  2   d_n = -0-1i 
assign u[4'b1110] [03] = 22'h 00001F;  // +0.1240334922877210 = 2^ 3 * ln( 1 +  0 * 2^(- 3+1) + ( 0^2+-1^2) * 2^(-2* 3) )   n =  3   d_n = -0-1i 
assign u[4'b1110] [04] = 22'h 00000F;  // +0.0623782466505195 = 2^ 4 * ln( 1 +  0 * 2^(- 4+1) + ( 0^2+-1^2) * 2^(-2* 4) )   n =  4   d_n = -0-1i 
assign u[4'b1110] [05] = 22'h 000007;  // +0.0312347511377731 = 2^ 5 * ln( 1 +  0 * 2^(- 5+1) + ( 0^2+-1^2) * 2^(-2* 5) )   n =  5   d_n = -0-1i 
assign u[4'b1110] [06] = 22'h 000003;  // +0.0156230929617406 = 2^ 6 * ln( 1 +  0 * 2^(- 6+1) + ( 0^2+-1^2) * 2^(-2* 6) )   n =  6   d_n = -0-1i 
assign u[4'b1110] [07] = 22'h 000001;  // +0.0078122615911219 = 2^ 7 * ln( 1 +  0 * 2^(- 7+1) + ( 0^2+-1^2) * 2^(-2* 7) )   n =  7   d_n = -0-1i 
assign u[4'b1110] [08] = 22'h 000000;  // +0.0039062201979808 = 2^ 8 * ln( 1 +  0 * 2^(- 8+1) + ( 0^2+-1^2) * 2^(-2* 8) )   n =  8   d_n = -0-1i 
assign u[4'b1110] [09] = 22'h 000000;  // +0.0019531212747156 = 2^ 9 * ln( 1 +  0 * 2^(- 9+1) + ( 0^2+-1^2) * 2^(-2* 9) )   n =  9   d_n = -0-1i 
assign u[4'b1110] [10] = 22'h 000000;  // +0.0009765620343389 = 2^10 * ln( 1 +  0 * 2^(-10+1) + ( 0^2+-1^2) * 2^(-2*10) )   n = 10   d_n = -0-1i 
assign u[4'b1110] [11] = 22'h 000000;  // +0.0004882811917923 = 2^11 * ln( 1 +  0 * 2^(-11+1) + ( 0^2+-1^2) * 2^(-2*11) )   n = 11   d_n = -0-1i 
assign u[4'b1110] [12] = 22'h 000000;  // +0.0002441406177240 = 2^12 * ln( 1 +  0 * 2^(-12+1) + ( 0^2+-1^2) * 2^(-2*12) )   n = 12   d_n = -0-1i 
assign u[4'b1110] [13] = 22'h 000000;  // +0.0001220703120453 = 2^13 * ln( 1 +  0 * 2^(-13+1) + ( 0^2+-1^2) * 2^(-2*13) )   n = 13   d_n = -0-1i 
assign u[4'b1110] [14] = 22'h 000000;  // +0.0000610351561932 = 2^14 * ln( 1 +  0 * 2^(-14+1) + ( 0^2+-1^2) * 2^(-2*14) )   n = 14   d_n = -0-1i 
assign u[4'b1110] [15] = 22'h 000000;  // +0.0000305175781179 = 2^15 * ln( 1 +  0 * 2^(-15+1) + ( 0^2+-1^2) * 2^(-2*15) )   n = 15   d_n = -0-1i 
assign u[4'b1110] [16] = 22'h 000000;  // +0.0000152587890616 = 2^16 * ln( 1 +  0 * 2^(-16+1) + ( 0^2+-1^2) * 2^(-2*16) )   n = 16   d_n = -0-1i 
assign u[4'b1110] [17] = 22'h 000000;  // +0.0000076293945311 = 2^17 * ln( 1 +  0 * 2^(-17+1) + ( 0^2+-1^2) * 2^(-2*17) )   n = 17   d_n = -0-1i 
assign u[4'b1110] [18] = 22'h 000000;  // +0.0000038146972656 = 2^18 * ln( 1 +  0 * 2^(-18+1) + ( 0^2+-1^2) * 2^(-2*18) )   n = 18   d_n = -0-1i 
assign u[4'b1110] [19] = 22'h 000000;  // +0.0000019073486328 = 2^19 * ln( 1 +  0 * 2^(-19+1) + ( 0^2+-1^2) * 2^(-2*19) )   n = 19   d_n = -0-1i 
assign u[4'b1110] [20] = 22'h 000000;  // +0.0000009536743164 = 2^20 * ln( 1 +  0 * 2^(-20+1) + ( 0^2+-1^2) * 2^(-2*20) )   n = 20   d_n = -0-1i 
assign u[4'b1110] [21] = 22'h 000000;  // +0.0000004768371582 = 2^21 * ln( 1 +  0 * 2^(-21+1) + ( 0^2+-1^2) * 2^(-2*21) )   n = 21   d_n = -0-1i 
assign u[4'b1110] [22] = 22'h 000000;  // +0.0000002384185791 = 2^22 * ln( 1 +  0 * 2^(-22+1) + ( 0^2+-1^2) * 2^(-2*22) )   n = 22   d_n = -0-1i 
assign u[4'b1110] [23] = 22'h 000000;  // +0.0000001192092896 = 2^23 * ln( 1 +  0 * 2^(-23+1) + ( 0^2+-1^2) * 2^(-2*23) )   n = 23   d_n = -0-1i 
assign u[4'b1110] [24] = 22'h 000000;  // +0.0000000596046448 = 2^24 * ln( 1 +  0 * 2^(-24+1) + ( 0^2+-1^2) * 2^(-2*24) )   n = 24   d_n = -0-1i 
assign u[4'b1110] [25] = 22'h 000000;  // +0.0000000298023224 = 2^25 * ln( 1 +  0 * 2^(-25+1) + ( 0^2+-1^2) * 2^(-2*25) )   n = 25   d_n = -0-1i 
assign u[4'b1110] [26] = 22'h 000000;  // +0.0000000000000000 = 2^26 * ln( 1 +  0 * 2^(-26+1) + ( 0^2+-1^2) * 2^(-2*26) )   n = 26   d_n = -0-1i 
assign u[4'b1110] [27] = 22'h 000000;  // +0.0000000000000000 = 2^27 * ln( 1 +  0 * 2^(-27+1) + ( 0^2+-1^2) * 2^(-2*27) )   n = 27   d_n = -0-1i 
assign u[4'b1110] [28] = 22'h 000000;  // +0.0000000000000000 = 2^28 * ln( 1 +  0 * 2^(-28+1) + ( 0^2+-1^2) * 2^(-2*28) )   n = 28   d_n = -0-1i 
assign u[4'b1110] [29] = 22'h 000000;  // +0.0000000000000000 = 2^29 * ln( 1 +  0 * 2^(-29+1) + ( 0^2+-1^2) * 2^(-2*29) )   n = 29   d_n = -0-1i 
assign u[4'b1110] [30] = 22'h 000000;  // +0.0000000000000000 = 2^30 * ln( 1 +  0 * 2^(-30+1) + ( 0^2+-1^2) * 2^(-2*30) )   n = 30   d_n = -0-1i 
assign u[4'b1110] [31] = 22'h 000000;  // +0.0000000000000000 = 2^31 * ln( 1 +  0 * 2^(-31+1) + ( 0^2+-1^2) * 2^(-2*31) )   n = 31   d_n = -0-1i 
assign u[4'b1110] [32] = 22'h 000000;  // +0.0000000000000000 = 2^32 * ln( 1 +  0 * 2^(-32+1) + ( 0^2+-1^2) * 2^(-2*32) )   n = 32   d_n = -0-1i 
assign u[4'b1110] [33] = 22'h 000000;  // +0.0000000000000000 = 2^33 * ln( 1 +  0 * 2^(-33+1) + ( 0^2+-1^2) * 2^(-2*33) )   n = 33   d_n = -0-1i 
assign u[4'b1110] [34] = 22'h 000000;  // +0.0000000000000000 = 2^34 * ln( 1 +  0 * 2^(-34+1) + ( 0^2+-1^2) * 2^(-2*34) )   n = 34   d_n = -0-1i 
assign u[4'b1110] [35] = 22'h 000000;  // +0.0000000000000000 = 2^35 * ln( 1 +  0 * 2^(-35+1) + ( 0^2+-1^2) * 2^(-2*35) )   n = 35   d_n = -0-1i 
assign u[4'b1110] [36] = 22'h 000000;  // +0.0000000000000000 = 2^36 * ln( 1 +  0 * 2^(-36+1) + ( 0^2+-1^2) * 2^(-2*36) )   n = 36   d_n = -0-1i 
assign u[4'b1110] [37] = 22'h 000000;  // +0.0000000000000000 = 2^37 * ln( 1 +  0 * 2^(-37+1) + ( 0^2+-1^2) * 2^(-2*37) )   n = 37   d_n = -0-1i 
assign u[4'b1110] [38] = 22'h 000000;  // +0.0000000000000000 = 2^38 * ln( 1 +  0 * 2^(-38+1) + ( 0^2+-1^2) * 2^(-2*38) )   n = 38   d_n = -0-1i 
assign u[4'b1110] [39] = 22'h 000000;  // +0.0000000000000000 = 2^39 * ln( 1 +  0 * 2^(-39+1) + ( 0^2+-1^2) * 2^(-2*39) )   n = 39   d_n = -0-1i 
assign u[4'b1110] [40] = 22'h 000000;  // +0.0000000000000000 = 2^40 * ln( 1 +  0 * 2^(-40+1) + ( 0^2+-1^2) * 2^(-2*40) )   n = 40   d_n = -0-1i 
assign u[4'b1110] [41] = 22'h 000000;  // +0.0000000000000000 = 2^41 * ln( 1 +  0 * 2^(-41+1) + ( 0^2+-1^2) * 2^(-2*41) )   n = 41   d_n = -0-1i 
assign u[4'b1110] [42] = 22'h 000000;  // +0.0000000000000000 = 2^42 * ln( 1 +  0 * 2^(-42+1) + ( 0^2+-1^2) * 2^(-2*42) )   n = 42   d_n = -0-1i 
assign u[4'b1110] [43] = 22'h 000000;  // +0.0000000000000000 = 2^43 * ln( 1 +  0 * 2^(-43+1) + ( 0^2+-1^2) * 2^(-2*43) )   n = 43   d_n = -0-1i 
assign u[4'b1110] [44] = 22'h 000000;  // +0.0000000000000000 = 2^44 * ln( 1 +  0 * 2^(-44+1) + ( 0^2+-1^2) * 2^(-2*44) )   n = 44   d_n = -0-1i 
assign u[4'b1110] [45] = 22'h 000000;  // +0.0000000000000000 = 2^45 * ln( 1 +  0 * 2^(-45+1) + ( 0^2+-1^2) * 2^(-2*45) )   n = 45   d_n = -0-1i 
assign u[4'b1110] [46] = 22'h 000000;  // +0.0000000000000000 = 2^46 * ln( 1 +  0 * 2^(-46+1) + ( 0^2+-1^2) * 2^(-2*46) )   n = 46   d_n = -0-1i 
assign u[4'b1110] [47] = 22'h 000000;  // +0.0000000000000000 = 2^47 * ln( 1 +  0 * 2^(-47+1) + ( 0^2+-1^2) * 2^(-2*47) )   n = 47   d_n = -0-1i 
assign u[4'b1110] [48] = 22'h 000000;  // +0.0000000000000000 = 2^48 * ln( 1 +  0 * 2^(-48+1) + ( 0^2+-1^2) * 2^(-2*48) )   n = 48   d_n = -0-1i 
assign u[4'b1110] [49] = 22'h 000000;  // +0.0000000000000000 = 2^49 * ln( 1 +  0 * 2^(-49+1) + ( 0^2+-1^2) * 2^(-2*49) )   n = 49   d_n = -0-1i 
assign u[4'b1110] [50] = 22'h 000000;  // +0.0000000000000000 = 2^50 * ln( 1 +  0 * 2^(-50+1) + ( 0^2+-1^2) * 2^(-2*50) )   n = 50   d_n = -0-1i 
assign u[4'b1110] [51] = 22'h 000000;  // +0.0000000000000000 = 2^51 * ln( 1 +  0 * 2^(-51+1) + ( 0^2+-1^2) * 2^(-2*51) )   n = 51   d_n = -0-1i 
assign u[4'b1110] [52] = 22'h 000000;  // +0.0000000000000000 = 2^52 * ln( 1 +  0 * 2^(-52+1) + ( 0^2+-1^2) * 2^(-2*52) )   n = 52   d_n = -0-1i 
assign u[4'b1110] [53] = 22'h 000000;  // +0.0000000000000000 = 2^53 * ln( 1 +  0 * 2^(-53+1) + ( 0^2+-1^2) * 2^(-2*53) )   n = 53   d_n = -0-1i 
assign u[4'b1110] [54] = 22'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 +  0 * 2^(-54+1) + ( 0^2+-1^2) * 2^(-2*54) )   n = 54   d_n = -0-1i 
assign u[4'b1110] [55] = 22'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 +  0 * 2^(-55+1) + ( 0^2+-1^2) * 2^(-2*55) )   n = 55   d_n = -0-1i 
assign u[4'b1110] [56] = 22'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 +  0 * 2^(-56+1) + ( 0^2+-1^2) * 2^(-2*56) )   n = 56   d_n = -0-1i 
assign u[4'b1110] [57] = 22'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 +  0 * 2^(-57+1) + ( 0^2+-1^2) * 2^(-2*57) )   n = 57   d_n = -0-1i 
assign u[4'b1110] [58] = 22'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 +  0 * 2^(-58+1) + ( 0^2+-1^2) * 2^(-2*58) )   n = 58   d_n = -0-1i 
assign u[4'b1110] [59] = 22'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 +  0 * 2^(-59+1) + ( 0^2+-1^2) * 2^(-2*59) )   n = 59   d_n = -0-1i 
assign u[4'b1110] [60] = 22'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 +  0 * 2^(-60+1) + ( 0^2+-1^2) * 2^(-2*60) )   n = 60   d_n = -0-1i 
assign u[4'b1110] [61] = 22'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 +  0 * 2^(-61+1) + ( 0^2+-1^2) * 2^(-2*61) )   n = 61   d_n = -0-1i 
assign u[4'b1110] [62] = 22'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 +  0 * 2^(-62+1) + ( 0^2+-1^2) * 2^(-2*62) )   n = 62   d_n = -0-1i 
assign u[4'b1110] [63] = 22'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 +  0 * 2^(-63+1) + ( 0^2+-1^2) * 2^(-2*63) )   n = 63   d_n = -0-1i 
assign u[4'b1110] [64] = 22'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 +  0 * 2^(-64+1) + ( 0^2+-1^2) * 2^(-2*64) )   n = 64   d_n = -0-1i 
assign u[4'b1111] [01] = 22'h 3FFE9D;  // -1.3862943611198904 = 2^ 1 * ln( 1 + -1 * 2^(- 1+1) + (-1^2+-1^2) * 2^(-2* 1) )   n =  1   d_n = -1-1i 
assign u[4'b1111] [02] = 22'h 3FFE1E;  // -1.8800145169829416 = 2^ 2 * ln( 1 + -1 * 2^(- 2+1) + (-1^2+-1^2) * 2^(-2* 2) )   n =  2   d_n = -1-1i 
assign u[4'b1111] [03] = 22'h 3FFE06;  // -1.9748806234522058 = 2^ 3 * ln( 1 + -1 * 2^(- 3+1) + (-1^2+-1^2) * 2^(-2* 3) )   n =  3   d_n = -1-1i 
assign u[4'b1111] [04] = 22'h 3FFE01;  // -1.9942791233164259 = 2^ 4 * ln( 1 + -1 * 2^(- 4+1) + (-1^2+-1^2) * 2^(-2* 4) )   n =  4   d_n = -1-1i 
assign u[4'b1111] [05] = 22'h 3FFE00;  // -1.9986353578798890 = 2^ 5 * ln( 1 + -1 * 2^(- 5+1) + (-1^2+-1^2) * 2^(-2* 5) )   n =  5   d_n = -1-1i 
assign u[4'b1111] [06] = 22'h 3FFE00;  // -1.9996667544388824 = 2^ 6 * ln( 1 + -1 * 2^(- 6+1) + (-1^2+-1^2) * 2^(-2* 6) )   n =  6   d_n = -1-1i 
assign u[4'b1111] [07] = 22'h 3FFE00;  // -1.9999176601574109 = 2^ 7 * ln( 1 + -1 * 2^(- 7+1) + (-1^2+-1^2) * 2^(-2* 7) )   n =  7   d_n = -1-1i 
assign u[4'b1111] [08] = 22'h 3FFE00;  // -1.9999795353661032 = 2^ 8 * ln( 1 + -1 * 2^(- 8+1) + (-1^2+-1^2) * 2^(-2* 8) )   n =  8   d_n = -1-1i 
assign u[4'b1111] [09] = 22'h 3FFE00;  // -1.9999948988125242 = 2^ 9 * ln( 1 + -1 * 2^(- 9+1) + (-1^2+-1^2) * 2^(-2* 9) )   n =  9   d_n = -1-1i 
assign u[4'b1111] [10] = 22'h 3FFE00;  // -1.9999987265701442 = 2^10 * ln( 1 + -1 * 2^(-10+1) + (-1^2+-1^2) * 2^(-2*10) )   n = 10   d_n = -1-1i 
assign u[4'b1111] [11] = 22'h 3FFE00;  // -1.9999996818756538 = 2^11 * ln( 1 + -1 * 2^(-11+1) + (-1^2+-1^2) * 2^(-2*11) )   n = 11   d_n = -1-1i 
assign u[4'b1111] [12] = 22'h 3FFE00;  // -1.9999999204980317 = 2^12 * ln( 1 + -1 * 2^(-12+1) + (-1^2+-1^2) * 2^(-2*12) )   n = 12   d_n = -1-1i 
assign u[4'b1111] [13] = 22'h 3FFE00;  // -1.9999999801276920 = 2^13 * ln( 1 + -1 * 2^(-13+1) + (-1^2+-1^2) * 2^(-2*13) )   n = 13   d_n = -1-1i 
assign u[4'b1111] [14] = 22'h 3FFE00;  // -1.9999999950326621 = 2^14 * ln( 1 + -1 * 2^(-14+1) + (-1^2+-1^2) * 2^(-2*14) )   n = 14   d_n = -1-1i 
assign u[4'b1111] [15] = 22'h 3FFE00;  // -1.9999999987582011 = 2^15 * ln( 1 + -1 * 2^(-15+1) + (-1^2+-1^2) * 2^(-2*15) )   n = 15   d_n = -1-1i 
assign u[4'b1111] [16] = 22'h 3FFE00;  // -1.9999999996895548 = 2^16 * ln( 1 + -1 * 2^(-16+1) + (-1^2+-1^2) * 2^(-2*16) )   n = 16   d_n = -1-1i 
assign u[4'b1111] [17] = 22'h 3FFE00;  // -1.9999999999223892 = 2^17 * ln( 1 + -1 * 2^(-17+1) + (-1^2+-1^2) * 2^(-2*17) )   n = 17   d_n = -1-1i 
assign u[4'b1111] [18] = 22'h 3FFE00;  // -1.9999999999951494 = 2^18 * ln( 1 + -1 * 2^(-18+1) + (-1^2+-1^2) * 2^(-2*18) )   n = 18   d_n = -1-1i 
assign u[4'b1111] [19] = 22'h 3FFE00;  // -1.9999999999987874 = 2^19 * ln( 1 + -1 * 2^(-19+1) + (-1^2+-1^2) * 2^(-2*19) )   n = 19   d_n = -1-1i 
assign u[4'b1111] [20] = 22'h 3FFE00;  // -1.9999999999996969 = 2^20 * ln( 1 + -1 * 2^(-20+1) + (-1^2+-1^2) * 2^(-2*20) )   n = 20   d_n = -1-1i 
assign u[4'b1111] [21] = 22'h 3FFE00;  // -1.9999999999999243 = 2^21 * ln( 1 + -1 * 2^(-21+1) + (-1^2+-1^2) * 2^(-2*21) )   n = 21   d_n = -1-1i 
assign u[4'b1111] [22] = 22'h 3FFE00;  // -1.9999999999999811 = 2^22 * ln( 1 + -1 * 2^(-22+1) + (-1^2+-1^2) * 2^(-2*22) )   n = 22   d_n = -1-1i 
assign u[4'b1111] [23] = 22'h 3FFE00;  // -1.9999999999999953 = 2^23 * ln( 1 + -1 * 2^(-23+1) + (-1^2+-1^2) * 2^(-2*23) )   n = 23   d_n = -1-1i 
assign u[4'b1111] [24] = 22'h 3FFE00;  // -1.9999999999999989 = 2^24 * ln( 1 + -1 * 2^(-24+1) + (-1^2+-1^2) * 2^(-2*24) )   n = 24   d_n = -1-1i 
assign u[4'b1111] [25] = 22'h 3FFE00;  // -1.9999999999999998 = 2^25 * ln( 1 + -1 * 2^(-25+1) + (-1^2+-1^2) * 2^(-2*25) )   n = 25   d_n = -1-1i 
assign u[4'b1111] [26] = 22'h 3FFE00;  // -2.0000000000000000 = 2^26 * ln( 1 + -1 * 2^(-26+1) + (-1^2+-1^2) * 2^(-2*26) )   n = 26   d_n = -1-1i 
assign u[4'b1111] [27] = 22'h 3FFDFF;  // -2.0000000074505806 = 2^27 * ln( 1 + -1 * 2^(-27+1) + (-1^2+-1^2) * 2^(-2*27) )   n = 27   d_n = -1-1i 
assign u[4'b1111] [28] = 22'h 3FFDFF;  // -2.0000000037252903 = 2^28 * ln( 1 + -1 * 2^(-28+1) + (-1^2+-1^2) * 2^(-2*28) )   n = 28   d_n = -1-1i 
assign u[4'b1111] [29] = 22'h 3FFDFF;  // -2.0000000018626451 = 2^29 * ln( 1 + -1 * 2^(-29+1) + (-1^2+-1^2) * 2^(-2*29) )   n = 29   d_n = -1-1i 
assign u[4'b1111] [30] = 22'h 3FFDFF;  // -2.0000000009313226 = 2^30 * ln( 1 + -1 * 2^(-30+1) + (-1^2+-1^2) * 2^(-2*30) )   n = 30   d_n = -1-1i 
assign u[4'b1111] [31] = 22'h 3FFDFF;  // -2.0000000004656613 = 2^31 * ln( 1 + -1 * 2^(-31+1) + (-1^2+-1^2) * 2^(-2*31) )   n = 31   d_n = -1-1i 
assign u[4'b1111] [32] = 22'h 3FFDFF;  // -2.0000000002328306 = 2^32 * ln( 1 + -1 * 2^(-32+1) + (-1^2+-1^2) * 2^(-2*32) )   n = 32   d_n = -1-1i 
assign u[4'b1111] [33] = 22'h 3FFDFF;  // -2.0000000001164153 = 2^33 * ln( 1 + -1 * 2^(-33+1) + (-1^2+-1^2) * 2^(-2*33) )   n = 33   d_n = -1-1i 
assign u[4'b1111] [34] = 22'h 3FFDFF;  // -2.0000000000582077 = 2^34 * ln( 1 + -1 * 2^(-34+1) + (-1^2+-1^2) * 2^(-2*34) )   n = 34   d_n = -1-1i 
assign u[4'b1111] [35] = 22'h 3FFDFF;  // -2.0000000000291038 = 2^35 * ln( 1 + -1 * 2^(-35+1) + (-1^2+-1^2) * 2^(-2*35) )   n = 35   d_n = -1-1i 
assign u[4'b1111] [36] = 22'h 3FFDFF;  // -2.0000000000145519 = 2^36 * ln( 1 + -1 * 2^(-36+1) + (-1^2+-1^2) * 2^(-2*36) )   n = 36   d_n = -1-1i 
assign u[4'b1111] [37] = 22'h 3FFDFF;  // -2.0000000000072760 = 2^37 * ln( 1 + -1 * 2^(-37+1) + (-1^2+-1^2) * 2^(-2*37) )   n = 37   d_n = -1-1i 
assign u[4'b1111] [38] = 22'h 3FFDFF;  // -2.0000000000036380 = 2^38 * ln( 1 + -1 * 2^(-38+1) + (-1^2+-1^2) * 2^(-2*38) )   n = 38   d_n = -1-1i 
assign u[4'b1111] [39] = 22'h 3FFDFF;  // -2.0000000000018190 = 2^39 * ln( 1 + -1 * 2^(-39+1) + (-1^2+-1^2) * 2^(-2*39) )   n = 39   d_n = -1-1i 
assign u[4'b1111] [40] = 22'h 3FFE00;  // -2.0000000000009095 = 2^40 * ln( 1 + -1 * 2^(-40+1) + (-1^2+-1^2) * 2^(-2*40) )   n = 40   d_n = -1-1i 
assign u[4'b1111] [41] = 22'h 3FFE00;  // -2.0000000000004547 = 2^41 * ln( 1 + -1 * 2^(-41+1) + (-1^2+-1^2) * 2^(-2*41) )   n = 41   d_n = -1-1i 
assign u[4'b1111] [42] = 22'h 3FFE00;  // -2.0000000000002274 = 2^42 * ln( 1 + -1 * 2^(-42+1) + (-1^2+-1^2) * 2^(-2*42) )   n = 42   d_n = -1-1i 
assign u[4'b1111] [43] = 22'h 3FFE00;  // -2.0000000000001137 = 2^43 * ln( 1 + -1 * 2^(-43+1) + (-1^2+-1^2) * 2^(-2*43) )   n = 43   d_n = -1-1i 
assign u[4'b1111] [44] = 22'h 3FFE00;  // -2.0000000000000568 = 2^44 * ln( 1 + -1 * 2^(-44+1) + (-1^2+-1^2) * 2^(-2*44) )   n = 44   d_n = -1-1i 
assign u[4'b1111] [45] = 22'h 3FFE00;  // -2.0000000000000284 = 2^45 * ln( 1 + -1 * 2^(-45+1) + (-1^2+-1^2) * 2^(-2*45) )   n = 45   d_n = -1-1i 
assign u[4'b1111] [46] = 22'h 3FFE00;  // -2.0000000000000142 = 2^46 * ln( 1 + -1 * 2^(-46+1) + (-1^2+-1^2) * 2^(-2*46) )   n = 46   d_n = -1-1i 
assign u[4'b1111] [47] = 22'h 3FFE00;  // -2.0000000000000071 = 2^47 * ln( 1 + -1 * 2^(-47+1) + (-1^2+-1^2) * 2^(-2*47) )   n = 47   d_n = -1-1i 
assign u[4'b1111] [48] = 22'h 3FFE00;  // -2.0000000000000036 = 2^48 * ln( 1 + -1 * 2^(-48+1) + (-1^2+-1^2) * 2^(-2*48) )   n = 48   d_n = -1-1i 
assign u[4'b1111] [49] = 22'h 3FFE00;  // -2.0000000000000018 = 2^49 * ln( 1 + -1 * 2^(-49+1) + (-1^2+-1^2) * 2^(-2*49) )   n = 49   d_n = -1-1i 
assign u[4'b1111] [50] = 22'h 3FFE00;  // -2.0000000000000009 = 2^50 * ln( 1 + -1 * 2^(-50+1) + (-1^2+-1^2) * 2^(-2*50) )   n = 50   d_n = -1-1i 
assign u[4'b1111] [51] = 22'h 3FFE00;  // -2.0000000000000004 = 2^51 * ln( 1 + -1 * 2^(-51+1) + (-1^2+-1^2) * 2^(-2*51) )   n = 51   d_n = -1-1i 
assign u[4'b1111] [52] = 22'h 3FFE00;  // -2.0000000000000004 = 2^52 * ln( 1 + -1 * 2^(-52+1) + (-1^2+-1^2) * 2^(-2*52) )   n = 52   d_n = -1-1i 
assign u[4'b1111] [53] = 22'h 3FFE00;  // -2.0000000000000000 = 2^53 * ln( 1 + -1 * 2^(-53+1) + (-1^2+-1^2) * 2^(-2*53) )   n = 53   d_n = -1-1i 
assign u[4'b1111] [54] = 22'h 000000;  // +0.0000000000000000 = 2^54 * ln( 1 + -1 * 2^(-54+1) + (-1^2+-1^2) * 2^(-2*54) )   n = 54   d_n = -1-1i 
assign u[4'b1111] [55] = 22'h 000000;  // +0.0000000000000000 = 2^55 * ln( 1 + -1 * 2^(-55+1) + (-1^2+-1^2) * 2^(-2*55) )   n = 55   d_n = -1-1i 
assign u[4'b1111] [56] = 22'h 000000;  // +0.0000000000000000 = 2^56 * ln( 1 + -1 * 2^(-56+1) + (-1^2+-1^2) * 2^(-2*56) )   n = 56   d_n = -1-1i 
assign u[4'b1111] [57] = 22'h 000000;  // +0.0000000000000000 = 2^57 * ln( 1 + -1 * 2^(-57+1) + (-1^2+-1^2) * 2^(-2*57) )   n = 57   d_n = -1-1i 
assign u[4'b1111] [58] = 22'h 000000;  // +0.0000000000000000 = 2^58 * ln( 1 + -1 * 2^(-58+1) + (-1^2+-1^2) * 2^(-2*58) )   n = 58   d_n = -1-1i 
assign u[4'b1111] [59] = 22'h 000000;  // +0.0000000000000000 = 2^59 * ln( 1 + -1 * 2^(-59+1) + (-1^2+-1^2) * 2^(-2*59) )   n = 59   d_n = -1-1i 
assign u[4'b1111] [60] = 22'h 000000;  // +0.0000000000000000 = 2^60 * ln( 1 + -1 * 2^(-60+1) + (-1^2+-1^2) * 2^(-2*60) )   n = 60   d_n = -1-1i 
assign u[4'b1111] [61] = 22'h 000000;  // +0.0000000000000000 = 2^61 * ln( 1 + -1 * 2^(-61+1) + (-1^2+-1^2) * 2^(-2*61) )   n = 61   d_n = -1-1i 
assign u[4'b1111] [62] = 22'h 000000;  // +0.0000000000000000 = 2^62 * ln( 1 + -1 * 2^(-62+1) + (-1^2+-1^2) * 2^(-2*62) )   n = 62   d_n = -1-1i 
assign u[4'b1111] [63] = 22'h 000000;  // +0.0000000000000000 = 2^63 * ln( 1 + -1 * 2^(-63+1) + (-1^2+-1^2) * 2^(-2*63) )   n = 63   d_n = -1-1i 
assign u[4'b1111] [64] = 22'h 000000;  // +0.0000000000000000 = 2^64 * ln( 1 + -1 * 2^(-64+1) + (-1^2+-1^2) * 2^(-2*64) )   n = 64   d_n = -1-1i 
assign v[4'b0000] [01] = 22'h 000000;  // +0.0000000000000000 = 2^(1+1) *  0 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = 0 
assign v[4'b0000] [02] = 22'h 000000;  // +0.0000000000000000 = 2^(2+1) *  0 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = 0 
assign v[4'b0000] [03] = 22'h 000000;  // +0.0000000000000000 = 2^(3+1) *  0 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = 0 
assign v[4'b0000] [04] = 22'h 000000;  // +0.0000000000000000 = 2^(4+1) *  0 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = 0 
assign v[4'b0000] [05] = 22'h 000000;  // +0.0000000000000000 = 2^(5+1) *  0 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = 0 
assign v[4'b0000] [06] = 22'h 000000;  // +0.0000000000000000 = 2^(6+1) *  0 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = 0 
assign v[4'b0000] [07] = 22'h 000000;  // +0.0000000000000000 = 2^(7+1) *  0 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = 0 
assign v[4'b0000] [08] = 22'h 000000;  // +0.0000000000000000 = 2^(8+1) *  0 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = 0 
assign v[4'b0000] [09] = 22'h 000000;  // +0.0000000000000000 = 2^(9+1) *  0 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = 0 
assign v[4'b0000] [10] = 22'h 000000;  // +0.0000000000000000 = 2^(10+1) *  0 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = 0 
assign v[4'b0000] [11] = 22'h 000000;  // +0.0000000000000000 = 2^(11+1) *  0 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = 0 
assign v[4'b0000] [12] = 22'h 000000;  // +0.0000000000000000 = 2^(12+1) *  0 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = 0 
assign v[4'b0000] [13] = 22'h 000000;  // +0.0000000000000000 = 2^(13+1) *  0 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = 0 
assign v[4'b0000] [14] = 22'h 000000;  // +0.0000000000000000 = 2^(14+1) *  0 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = 0 
assign v[4'b0000] [15] = 22'h 000000;  // +0.0000000000000000 = 2^(15+1) *  0 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = 0 
assign v[4'b0000] [16] = 22'h 000000;  // +0.0000000000000000 = 2^(16+1) *  0 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = 0 
assign v[4'b0000] [17] = 22'h 000000;  // +0.0000000000000000 = 2^(17+1) *  0 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = 0 
assign v[4'b0000] [18] = 22'h 000000;  // +0.0000000000000000 = 2^(18+1) *  0 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = 0 
assign v[4'b0000] [19] = 22'h 000000;  // +0.0000000000000000 = 2^(19+1) *  0 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = 0 
assign v[4'b0000] [20] = 22'h 000000;  // +0.0000000000000000 = 2^(20+1) *  0 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = 0 
assign v[4'b0000] [21] = 22'h 000000;  // +0.0000000000000000 = 2^(21+1) *  0 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = 0 
assign v[4'b0000] [22] = 22'h 000000;  // +0.0000000000000000 = 2^(22+1) *  0 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = 0 
assign v[4'b0000] [23] = 22'h 000000;  // +0.0000000000000000 = 2^(23+1) *  0 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = 0 
assign v[4'b0000] [24] = 22'h 000000;  // +0.0000000000000000 = 2^(24+1) *  0 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = 0 
assign v[4'b0000] [25] = 22'h 000000;  // +0.0000000000000000 = 2^(25+1) *  0 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = 0 
assign v[4'b0000] [26] = 22'h 000000;  // +0.0000000000000000 = 2^(26+1) *  0 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = 0 
assign v[4'b0000] [27] = 22'h 000000;  // +0.0000000000000000 = 2^(27+1) *  0 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = 0 
assign v[4'b0000] [28] = 22'h 000000;  // +0.0000000000000000 = 2^(28+1) *  0 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = 0 
assign v[4'b0000] [29] = 22'h 000000;  // +0.0000000000000000 = 2^(29+1) *  0 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = 0 
assign v[4'b0000] [30] = 22'h 000000;  // +0.0000000000000000 = 2^(30+1) *  0 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = 0 
assign v[4'b0000] [31] = 22'h 000000;  // +0.0000000000000000 = 2^(31+1) *  0 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = 0 
assign v[4'b0000] [32] = 22'h 000000;  // +0.0000000000000000 = 2^(32+1) *  0 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = 0 
assign v[4'b0000] [33] = 22'h 000000;  // +0.0000000000000000 = 2^(33+1) *  0 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = 0 
assign v[4'b0000] [34] = 22'h 000000;  // +0.0000000000000000 = 2^(34+1) *  0 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = 0 
assign v[4'b0000] [35] = 22'h 000000;  // +0.0000000000000000 = 2^(35+1) *  0 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = 0 
assign v[4'b0000] [36] = 22'h 000000;  // +0.0000000000000000 = 2^(36+1) *  0 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = 0 
assign v[4'b0000] [37] = 22'h 000000;  // +0.0000000000000000 = 2^(37+1) *  0 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = 0 
assign v[4'b0000] [38] = 22'h 000000;  // +0.0000000000000000 = 2^(38+1) *  0 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = 0 
assign v[4'b0000] [39] = 22'h 000000;  // +0.0000000000000000 = 2^(39+1) *  0 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = 0 
assign v[4'b0000] [40] = 22'h 000000;  // +0.0000000000000000 = 2^(40+1) *  0 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = 0 
assign v[4'b0000] [41] = 22'h 000000;  // +0.0000000000000000 = 2^(41+1) *  0 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = 0 
assign v[4'b0000] [42] = 22'h 000000;  // +0.0000000000000000 = 2^(42+1) *  0 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = 0 
assign v[4'b0000] [43] = 22'h 000000;  // +0.0000000000000000 = 2^(43+1) *  0 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = 0 
assign v[4'b0000] [44] = 22'h 000000;  // +0.0000000000000000 = 2^(44+1) *  0 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = 0 
assign v[4'b0000] [45] = 22'h 000000;  // +0.0000000000000000 = 2^(45+1) *  0 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = 0 
assign v[4'b0000] [46] = 22'h 000000;  // +0.0000000000000000 = 2^(46+1) *  0 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = 0 
assign v[4'b0000] [47] = 22'h 000000;  // +0.0000000000000000 = 2^(47+1) *  0 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = 0 
assign v[4'b0000] [48] = 22'h 000000;  // +0.0000000000000000 = 2^(48+1) *  0 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = 0 
assign v[4'b0000] [49] = 22'h 000000;  // +0.0000000000000000 = 2^(49+1) *  0 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = 0 
assign v[4'b0000] [50] = 22'h 000000;  // +0.0000000000000000 = 2^(50+1) *  0 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = 0 
assign v[4'b0000] [51] = 22'h 000000;  // +0.0000000000000000 = 2^(51+1) *  0 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = 0 
assign v[4'b0000] [52] = 22'h 000000;  // +0.0000000000000000 = 2^(52+1) *  0 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = 0 
assign v[4'b0000] [53] = 22'h 000000;  // +0.0000000000000000 = 2^(53+1) *  0 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = 0 
assign v[4'b0000] [54] = 22'h 000000;  // +0.0000000000000000 = 2^(54+1) *  0 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = 0 
assign v[4'b0000] [55] = 22'h 000000;  // +0.0000000000000000 = 2^(55+1) *  0 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = 0 
assign v[4'b0000] [56] = 22'h 000000;  // +0.0000000000000000 = 2^(56+1) *  0 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = 0 
assign v[4'b0000] [57] = 22'h 000000;  // +0.0000000000000000 = 2^(57+1) *  0 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = 0 
assign v[4'b0000] [58] = 22'h 000000;  // +0.0000000000000000 = 2^(58+1) *  0 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = 0 
assign v[4'b0000] [59] = 22'h 000000;  // +0.0000000000000000 = 2^(59+1) *  0 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = 0 
assign v[4'b0000] [60] = 22'h 000000;  // +0.0000000000000000 = 2^(60+1) *  0 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = 0 
assign v[4'b0000] [61] = 22'h 000000;  // +0.0000000000000000 = 2^(61+1) *  0 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = 0 
assign v[4'b0000] [62] = 22'h 000000;  // +0.0000000000000000 = 2^(62+1) *  0 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = 0 
assign v[4'b0000] [63] = 22'h 000000;  // +0.0000000000000000 = 2^(63+1) *  0 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = 0 
assign v[4'b0000] [64] = 22'h 000000;  // +0.0000000000000000 = 2^(64+1) *  0 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = 0 
assign v[4'b0001] [01] = 22'h 000000;  // +0.0000000000000000 = 2^(1+1) *  0 * atan( 1 / (  1 + 2^1 ) )   n =  1   d_n = 1 
assign v[4'b0001] [02] = 22'h 000000;  // +0.0000000000000000 = 2^(2+1) *  0 * atan( 1 / (  1 + 2^2 ) )   n =  2   d_n = 1 
assign v[4'b0001] [03] = 22'h 000000;  // +0.0000000000000000 = 2^(3+1) *  0 * atan( 1 / (  1 + 2^3 ) )   n =  3   d_n = 1 
assign v[4'b0001] [04] = 22'h 000000;  // +0.0000000000000000 = 2^(4+1) *  0 * atan( 1 / (  1 + 2^4 ) )   n =  4   d_n = 1 
assign v[4'b0001] [05] = 22'h 000000;  // +0.0000000000000000 = 2^(5+1) *  0 * atan( 1 / (  1 + 2^5 ) )   n =  5   d_n = 1 
assign v[4'b0001] [06] = 22'h 000000;  // +0.0000000000000000 = 2^(6+1) *  0 * atan( 1 / (  1 + 2^6 ) )   n =  6   d_n = 1 
assign v[4'b0001] [07] = 22'h 000000;  // +0.0000000000000000 = 2^(7+1) *  0 * atan( 1 / (  1 + 2^7 ) )   n =  7   d_n = 1 
assign v[4'b0001] [08] = 22'h 000000;  // +0.0000000000000000 = 2^(8+1) *  0 * atan( 1 / (  1 + 2^8 ) )   n =  8   d_n = 1 
assign v[4'b0001] [09] = 22'h 000000;  // +0.0000000000000000 = 2^(9+1) *  0 * atan( 1 / (  1 + 2^9 ) )   n =  9   d_n = 1 
assign v[4'b0001] [10] = 22'h 000000;  // +0.0000000000000000 = 2^(10+1) *  0 * atan( 1 / (  1 + 2^10 ) )   n = 10   d_n = 1 
assign v[4'b0001] [11] = 22'h 000000;  // +0.0000000000000000 = 2^(11+1) *  0 * atan( 1 / (  1 + 2^11 ) )   n = 11   d_n = 1 
assign v[4'b0001] [12] = 22'h 000000;  // +0.0000000000000000 = 2^(12+1) *  0 * atan( 1 / (  1 + 2^12 ) )   n = 12   d_n = 1 
assign v[4'b0001] [13] = 22'h 000000;  // +0.0000000000000000 = 2^(13+1) *  0 * atan( 1 / (  1 + 2^13 ) )   n = 13   d_n = 1 
assign v[4'b0001] [14] = 22'h 000000;  // +0.0000000000000000 = 2^(14+1) *  0 * atan( 1 / (  1 + 2^14 ) )   n = 14   d_n = 1 
assign v[4'b0001] [15] = 22'h 000000;  // +0.0000000000000000 = 2^(15+1) *  0 * atan( 1 / (  1 + 2^15 ) )   n = 15   d_n = 1 
assign v[4'b0001] [16] = 22'h 000000;  // +0.0000000000000000 = 2^(16+1) *  0 * atan( 1 / (  1 + 2^16 ) )   n = 16   d_n = 1 
assign v[4'b0001] [17] = 22'h 000000;  // +0.0000000000000000 = 2^(17+1) *  0 * atan( 1 / (  1 + 2^17 ) )   n = 17   d_n = 1 
assign v[4'b0001] [18] = 22'h 000000;  // +0.0000000000000000 = 2^(18+1) *  0 * atan( 1 / (  1 + 2^18 ) )   n = 18   d_n = 1 
assign v[4'b0001] [19] = 22'h 000000;  // +0.0000000000000000 = 2^(19+1) *  0 * atan( 1 / (  1 + 2^19 ) )   n = 19   d_n = 1 
assign v[4'b0001] [20] = 22'h 000000;  // +0.0000000000000000 = 2^(20+1) *  0 * atan( 1 / (  1 + 2^20 ) )   n = 20   d_n = 1 
assign v[4'b0001] [21] = 22'h 000000;  // +0.0000000000000000 = 2^(21+1) *  0 * atan( 1 / (  1 + 2^21 ) )   n = 21   d_n = 1 
assign v[4'b0001] [22] = 22'h 000000;  // +0.0000000000000000 = 2^(22+1) *  0 * atan( 1 / (  1 + 2^22 ) )   n = 22   d_n = 1 
assign v[4'b0001] [23] = 22'h 000000;  // +0.0000000000000000 = 2^(23+1) *  0 * atan( 1 / (  1 + 2^23 ) )   n = 23   d_n = 1 
assign v[4'b0001] [24] = 22'h 000000;  // +0.0000000000000000 = 2^(24+1) *  0 * atan( 1 / (  1 + 2^24 ) )   n = 24   d_n = 1 
assign v[4'b0001] [25] = 22'h 000000;  // +0.0000000000000000 = 2^(25+1) *  0 * atan( 1 / (  1 + 2^25 ) )   n = 25   d_n = 1 
assign v[4'b0001] [26] = 22'h 000000;  // +0.0000000000000000 = 2^(26+1) *  0 * atan( 1 / (  1 + 2^26 ) )   n = 26   d_n = 1 
assign v[4'b0001] [27] = 22'h 000000;  // +0.0000000000000000 = 2^(27+1) *  0 * atan( 1 / (  1 + 2^27 ) )   n = 27   d_n = 1 
assign v[4'b0001] [28] = 22'h 000000;  // +0.0000000000000000 = 2^(28+1) *  0 * atan( 1 / (  1 + 2^28 ) )   n = 28   d_n = 1 
assign v[4'b0001] [29] = 22'h 000000;  // +0.0000000000000000 = 2^(29+1) *  0 * atan( 1 / (  1 + 2^29 ) )   n = 29   d_n = 1 
assign v[4'b0001] [30] = 22'h 000000;  // +0.0000000000000000 = 2^(30+1) *  0 * atan( 1 / (  1 + 2^30 ) )   n = 30   d_n = 1 
assign v[4'b0001] [31] = 22'h 000000;  // +0.0000000000000000 = 2^(31+1) *  0 * atan( 1 / (  1 + 2^31 ) )   n = 31   d_n = 1 
assign v[4'b0001] [32] = 22'h 000000;  // +0.0000000000000000 = 2^(32+1) *  0 * atan( 1 / (  1 + 2^32 ) )   n = 32   d_n = 1 
assign v[4'b0001] [33] = 22'h 000000;  // +0.0000000000000000 = 2^(33+1) *  0 * atan( 1 / (  1 + 2^33 ) )   n = 33   d_n = 1 
assign v[4'b0001] [34] = 22'h 000000;  // +0.0000000000000000 = 2^(34+1) *  0 * atan( 1 / (  1 + 2^34 ) )   n = 34   d_n = 1 
assign v[4'b0001] [35] = 22'h 000000;  // +0.0000000000000000 = 2^(35+1) *  0 * atan( 1 / (  1 + 2^35 ) )   n = 35   d_n = 1 
assign v[4'b0001] [36] = 22'h 000000;  // +0.0000000000000000 = 2^(36+1) *  0 * atan( 1 / (  1 + 2^36 ) )   n = 36   d_n = 1 
assign v[4'b0001] [37] = 22'h 000000;  // +0.0000000000000000 = 2^(37+1) *  0 * atan( 1 / (  1 + 2^37 ) )   n = 37   d_n = 1 
assign v[4'b0001] [38] = 22'h 000000;  // +0.0000000000000000 = 2^(38+1) *  0 * atan( 1 / (  1 + 2^38 ) )   n = 38   d_n = 1 
assign v[4'b0001] [39] = 22'h 000000;  // +0.0000000000000000 = 2^(39+1) *  0 * atan( 1 / (  1 + 2^39 ) )   n = 39   d_n = 1 
assign v[4'b0001] [40] = 22'h 000000;  // +0.0000000000000000 = 2^(40+1) *  0 * atan( 1 / (  1 + 2^40 ) )   n = 40   d_n = 1 
assign v[4'b0001] [41] = 22'h 000000;  // +0.0000000000000000 = 2^(41+1) *  0 * atan( 1 / (  1 + 2^41 ) )   n = 41   d_n = 1 
assign v[4'b0001] [42] = 22'h 000000;  // +0.0000000000000000 = 2^(42+1) *  0 * atan( 1 / (  1 + 2^42 ) )   n = 42   d_n = 1 
assign v[4'b0001] [43] = 22'h 000000;  // +0.0000000000000000 = 2^(43+1) *  0 * atan( 1 / (  1 + 2^43 ) )   n = 43   d_n = 1 
assign v[4'b0001] [44] = 22'h 000000;  // +0.0000000000000000 = 2^(44+1) *  0 * atan( 1 / (  1 + 2^44 ) )   n = 44   d_n = 1 
assign v[4'b0001] [45] = 22'h 000000;  // +0.0000000000000000 = 2^(45+1) *  0 * atan( 1 / (  1 + 2^45 ) )   n = 45   d_n = 1 
assign v[4'b0001] [46] = 22'h 000000;  // +0.0000000000000000 = 2^(46+1) *  0 * atan( 1 / (  1 + 2^46 ) )   n = 46   d_n = 1 
assign v[4'b0001] [47] = 22'h 000000;  // +0.0000000000000000 = 2^(47+1) *  0 * atan( 1 / (  1 + 2^47 ) )   n = 47   d_n = 1 
assign v[4'b0001] [48] = 22'h 000000;  // +0.0000000000000000 = 2^(48+1) *  0 * atan( 1 / (  1 + 2^48 ) )   n = 48   d_n = 1 
assign v[4'b0001] [49] = 22'h 000000;  // +0.0000000000000000 = 2^(49+1) *  0 * atan( 1 / (  1 + 2^49 ) )   n = 49   d_n = 1 
assign v[4'b0001] [50] = 22'h 000000;  // +0.0000000000000000 = 2^(50+1) *  0 * atan( 1 / (  1 + 2^50 ) )   n = 50   d_n = 1 
assign v[4'b0001] [51] = 22'h 000000;  // +0.0000000000000000 = 2^(51+1) *  0 * atan( 1 / (  1 + 2^51 ) )   n = 51   d_n = 1 
assign v[4'b0001] [52] = 22'h 000000;  // +0.0000000000000000 = 2^(52+1) *  0 * atan( 1 / (  1 + 2^52 ) )   n = 52   d_n = 1 
assign v[4'b0001] [53] = 22'h 000000;  // +0.0000000000000000 = 2^(53+1) *  0 * atan( 1 / (  1 + 2^53 ) )   n = 53   d_n = 1 
assign v[4'b0001] [54] = 22'h 000000;  // +0.0000000000000000 = 2^(54+1) *  0 * atan( 1 / (  1 + 2^54 ) )   n = 54   d_n = 1 
assign v[4'b0001] [55] = 22'h 000000;  // +0.0000000000000000 = 2^(55+1) *  0 * atan( 1 / (  1 + 2^55 ) )   n = 55   d_n = 1 
assign v[4'b0001] [56] = 22'h 000000;  // +0.0000000000000000 = 2^(56+1) *  0 * atan( 1 / (  1 + 2^56 ) )   n = 56   d_n = 1 
assign v[4'b0001] [57] = 22'h 000000;  // +0.0000000000000000 = 2^(57+1) *  0 * atan( 1 / (  1 + 2^57 ) )   n = 57   d_n = 1 
assign v[4'b0001] [58] = 22'h 000000;  // +0.0000000000000000 = 2^(58+1) *  0 * atan( 1 / (  1 + 2^58 ) )   n = 58   d_n = 1 
assign v[4'b0001] [59] = 22'h 000000;  // +0.0000000000000000 = 2^(59+1) *  0 * atan( 1 / (  1 + 2^59 ) )   n = 59   d_n = 1 
assign v[4'b0001] [60] = 22'h 000000;  // +0.0000000000000000 = 2^(60+1) *  0 * atan( 1 / (  1 + 2^60 ) )   n = 60   d_n = 1 
assign v[4'b0001] [61] = 22'h 000000;  // +0.0000000000000000 = 2^(61+1) *  0 * atan( 1 / (  1 + 2^61 ) )   n = 61   d_n = 1 
assign v[4'b0001] [62] = 22'h 000000;  // +0.0000000000000000 = 2^(62+1) *  0 * atan( 1 / (  1 + 2^62 ) )   n = 62   d_n = 1 
assign v[4'b0001] [63] = 22'h 000000;  // +0.0000000000000000 = 2^(63+1) *  0 * atan( 1 / (  1 + 2^63 ) )   n = 63   d_n = 1 
assign v[4'b0001] [64] = 22'h 000000;  // +0.0000000000000000 = 2^(64+1) *  0 * atan( 1 / (  1 + 2^64 ) )   n = 64   d_n = 1 
assign v[4'b0010] [01] = 22'h 000000;  // +0.0000000000000000 = 2^(1+1) *  0 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = -0 
assign v[4'b0010] [02] = 22'h 000000;  // +0.0000000000000000 = 2^(2+1) *  0 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = -0 
assign v[4'b0010] [03] = 22'h 000000;  // +0.0000000000000000 = 2^(3+1) *  0 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = -0 
assign v[4'b0010] [04] = 22'h 000000;  // +0.0000000000000000 = 2^(4+1) *  0 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = -0 
assign v[4'b0010] [05] = 22'h 000000;  // +0.0000000000000000 = 2^(5+1) *  0 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = -0 
assign v[4'b0010] [06] = 22'h 000000;  // +0.0000000000000000 = 2^(6+1) *  0 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = -0 
assign v[4'b0010] [07] = 22'h 000000;  // +0.0000000000000000 = 2^(7+1) *  0 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = -0 
assign v[4'b0010] [08] = 22'h 000000;  // +0.0000000000000000 = 2^(8+1) *  0 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = -0 
assign v[4'b0010] [09] = 22'h 000000;  // +0.0000000000000000 = 2^(9+1) *  0 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = -0 
assign v[4'b0010] [10] = 22'h 000000;  // +0.0000000000000000 = 2^(10+1) *  0 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = -0 
assign v[4'b0010] [11] = 22'h 000000;  // +0.0000000000000000 = 2^(11+1) *  0 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = -0 
assign v[4'b0010] [12] = 22'h 000000;  // +0.0000000000000000 = 2^(12+1) *  0 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = -0 
assign v[4'b0010] [13] = 22'h 000000;  // +0.0000000000000000 = 2^(13+1) *  0 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = -0 
assign v[4'b0010] [14] = 22'h 000000;  // +0.0000000000000000 = 2^(14+1) *  0 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = -0 
assign v[4'b0010] [15] = 22'h 000000;  // +0.0000000000000000 = 2^(15+1) *  0 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = -0 
assign v[4'b0010] [16] = 22'h 000000;  // +0.0000000000000000 = 2^(16+1) *  0 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = -0 
assign v[4'b0010] [17] = 22'h 000000;  // +0.0000000000000000 = 2^(17+1) *  0 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = -0 
assign v[4'b0010] [18] = 22'h 000000;  // +0.0000000000000000 = 2^(18+1) *  0 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = -0 
assign v[4'b0010] [19] = 22'h 000000;  // +0.0000000000000000 = 2^(19+1) *  0 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = -0 
assign v[4'b0010] [20] = 22'h 000000;  // +0.0000000000000000 = 2^(20+1) *  0 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = -0 
assign v[4'b0010] [21] = 22'h 000000;  // +0.0000000000000000 = 2^(21+1) *  0 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = -0 
assign v[4'b0010] [22] = 22'h 000000;  // +0.0000000000000000 = 2^(22+1) *  0 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = -0 
assign v[4'b0010] [23] = 22'h 000000;  // +0.0000000000000000 = 2^(23+1) *  0 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = -0 
assign v[4'b0010] [24] = 22'h 000000;  // +0.0000000000000000 = 2^(24+1) *  0 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = -0 
assign v[4'b0010] [25] = 22'h 000000;  // +0.0000000000000000 = 2^(25+1) *  0 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = -0 
assign v[4'b0010] [26] = 22'h 000000;  // +0.0000000000000000 = 2^(26+1) *  0 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = -0 
assign v[4'b0010] [27] = 22'h 000000;  // +0.0000000000000000 = 2^(27+1) *  0 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = -0 
assign v[4'b0010] [28] = 22'h 000000;  // +0.0000000000000000 = 2^(28+1) *  0 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = -0 
assign v[4'b0010] [29] = 22'h 000000;  // +0.0000000000000000 = 2^(29+1) *  0 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = -0 
assign v[4'b0010] [30] = 22'h 000000;  // +0.0000000000000000 = 2^(30+1) *  0 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = -0 
assign v[4'b0010] [31] = 22'h 000000;  // +0.0000000000000000 = 2^(31+1) *  0 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = -0 
assign v[4'b0010] [32] = 22'h 000000;  // +0.0000000000000000 = 2^(32+1) *  0 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = -0 
assign v[4'b0010] [33] = 22'h 000000;  // +0.0000000000000000 = 2^(33+1) *  0 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = -0 
assign v[4'b0010] [34] = 22'h 000000;  // +0.0000000000000000 = 2^(34+1) *  0 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = -0 
assign v[4'b0010] [35] = 22'h 000000;  // +0.0000000000000000 = 2^(35+1) *  0 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = -0 
assign v[4'b0010] [36] = 22'h 000000;  // +0.0000000000000000 = 2^(36+1) *  0 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = -0 
assign v[4'b0010] [37] = 22'h 000000;  // +0.0000000000000000 = 2^(37+1) *  0 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = -0 
assign v[4'b0010] [38] = 22'h 000000;  // +0.0000000000000000 = 2^(38+1) *  0 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = -0 
assign v[4'b0010] [39] = 22'h 000000;  // +0.0000000000000000 = 2^(39+1) *  0 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = -0 
assign v[4'b0010] [40] = 22'h 000000;  // +0.0000000000000000 = 2^(40+1) *  0 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = -0 
assign v[4'b0010] [41] = 22'h 000000;  // +0.0000000000000000 = 2^(41+1) *  0 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = -0 
assign v[4'b0010] [42] = 22'h 000000;  // +0.0000000000000000 = 2^(42+1) *  0 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = -0 
assign v[4'b0010] [43] = 22'h 000000;  // +0.0000000000000000 = 2^(43+1) *  0 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = -0 
assign v[4'b0010] [44] = 22'h 000000;  // +0.0000000000000000 = 2^(44+1) *  0 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = -0 
assign v[4'b0010] [45] = 22'h 000000;  // +0.0000000000000000 = 2^(45+1) *  0 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = -0 
assign v[4'b0010] [46] = 22'h 000000;  // +0.0000000000000000 = 2^(46+1) *  0 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = -0 
assign v[4'b0010] [47] = 22'h 000000;  // +0.0000000000000000 = 2^(47+1) *  0 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = -0 
assign v[4'b0010] [48] = 22'h 000000;  // +0.0000000000000000 = 2^(48+1) *  0 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = -0 
assign v[4'b0010] [49] = 22'h 000000;  // +0.0000000000000000 = 2^(49+1) *  0 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = -0 
assign v[4'b0010] [50] = 22'h 000000;  // +0.0000000000000000 = 2^(50+1) *  0 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = -0 
assign v[4'b0010] [51] = 22'h 000000;  // +0.0000000000000000 = 2^(51+1) *  0 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = -0 
assign v[4'b0010] [52] = 22'h 000000;  // +0.0000000000000000 = 2^(52+1) *  0 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = -0 
assign v[4'b0010] [53] = 22'h 000000;  // +0.0000000000000000 = 2^(53+1) *  0 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = -0 
assign v[4'b0010] [54] = 22'h 000000;  // +0.0000000000000000 = 2^(54+1) *  0 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = -0 
assign v[4'b0010] [55] = 22'h 000000;  // +0.0000000000000000 = 2^(55+1) *  0 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = -0 
assign v[4'b0010] [56] = 22'h 000000;  // +0.0000000000000000 = 2^(56+1) *  0 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = -0 
assign v[4'b0010] [57] = 22'h 000000;  // +0.0000000000000000 = 2^(57+1) *  0 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = -0 
assign v[4'b0010] [58] = 22'h 000000;  // +0.0000000000000000 = 2^(58+1) *  0 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = -0 
assign v[4'b0010] [59] = 22'h 000000;  // +0.0000000000000000 = 2^(59+1) *  0 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = -0 
assign v[4'b0010] [60] = 22'h 000000;  // +0.0000000000000000 = 2^(60+1) *  0 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = -0 
assign v[4'b0010] [61] = 22'h 000000;  // +0.0000000000000000 = 2^(61+1) *  0 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = -0 
assign v[4'b0010] [62] = 22'h 000000;  // +0.0000000000000000 = 2^(62+1) *  0 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = -0 
assign v[4'b0010] [63] = 22'h 000000;  // +0.0000000000000000 = 2^(63+1) *  0 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = -0 
assign v[4'b0010] [64] = 22'h 000000;  // +0.0000000000000000 = 2^(64+1) *  0 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = -0 
assign v[4'b0011] [01] = 22'h 000000;  // -0.0000000000000000 = 2^(1+1) *  0 * atan( 1 / ( -1 + 2^1 ) )   n =  1   d_n = -1 
assign v[4'b0011] [02] = 22'h 000000;  // -0.0000000000000000 = 2^(2+1) *  0 * atan( 1 / ( -1 + 2^2 ) )   n =  2   d_n = -1 
assign v[4'b0011] [03] = 22'h 000000;  // -0.0000000000000000 = 2^(3+1) *  0 * atan( 1 / ( -1 + 2^3 ) )   n =  3   d_n = -1 
assign v[4'b0011] [04] = 22'h 000000;  // -0.0000000000000000 = 2^(4+1) *  0 * atan( 1 / ( -1 + 2^4 ) )   n =  4   d_n = -1 
assign v[4'b0011] [05] = 22'h 000000;  // -0.0000000000000000 = 2^(5+1) *  0 * atan( 1 / ( -1 + 2^5 ) )   n =  5   d_n = -1 
assign v[4'b0011] [06] = 22'h 000000;  // -0.0000000000000000 = 2^(6+1) *  0 * atan( 1 / ( -1 + 2^6 ) )   n =  6   d_n = -1 
assign v[4'b0011] [07] = 22'h 000000;  // -0.0000000000000000 = 2^(7+1) *  0 * atan( 1 / ( -1 + 2^7 ) )   n =  7   d_n = -1 
assign v[4'b0011] [08] = 22'h 000000;  // -0.0000000000000000 = 2^(8+1) *  0 * atan( 1 / ( -1 + 2^8 ) )   n =  8   d_n = -1 
assign v[4'b0011] [09] = 22'h 000000;  // -0.0000000000000000 = 2^(9+1) *  0 * atan( 1 / ( -1 + 2^9 ) )   n =  9   d_n = -1 
assign v[4'b0011] [10] = 22'h 000000;  // -0.0000000000000000 = 2^(10+1) *  0 * atan( 1 / ( -1 + 2^10 ) )   n = 10   d_n = -1 
assign v[4'b0011] [11] = 22'h 000000;  // -0.0000000000000000 = 2^(11+1) *  0 * atan( 1 / ( -1 + 2^11 ) )   n = 11   d_n = -1 
assign v[4'b0011] [12] = 22'h 000000;  // -0.0000000000000000 = 2^(12+1) *  0 * atan( 1 / ( -1 + 2^12 ) )   n = 12   d_n = -1 
assign v[4'b0011] [13] = 22'h 000000;  // -0.0000000000000000 = 2^(13+1) *  0 * atan( 1 / ( -1 + 2^13 ) )   n = 13   d_n = -1 
assign v[4'b0011] [14] = 22'h 000000;  // -0.0000000000000000 = 2^(14+1) *  0 * atan( 1 / ( -1 + 2^14 ) )   n = 14   d_n = -1 
assign v[4'b0011] [15] = 22'h 000000;  // -0.0000000000000000 = 2^(15+1) *  0 * atan( 1 / ( -1 + 2^15 ) )   n = 15   d_n = -1 
assign v[4'b0011] [16] = 22'h 000000;  // -0.0000000000000000 = 2^(16+1) *  0 * atan( 1 / ( -1 + 2^16 ) )   n = 16   d_n = -1 
assign v[4'b0011] [17] = 22'h 000000;  // -0.0000000000000000 = 2^(17+1) *  0 * atan( 1 / ( -1 + 2^17 ) )   n = 17   d_n = -1 
assign v[4'b0011] [18] = 22'h 000000;  // -0.0000000000000000 = 2^(18+1) *  0 * atan( 1 / ( -1 + 2^18 ) )   n = 18   d_n = -1 
assign v[4'b0011] [19] = 22'h 000000;  // -0.0000000000000000 = 2^(19+1) *  0 * atan( 1 / ( -1 + 2^19 ) )   n = 19   d_n = -1 
assign v[4'b0011] [20] = 22'h 000000;  // -0.0000000000000000 = 2^(20+1) *  0 * atan( 1 / ( -1 + 2^20 ) )   n = 20   d_n = -1 
assign v[4'b0011] [21] = 22'h 000000;  // -0.0000000000000000 = 2^(21+1) *  0 * atan( 1 / ( -1 + 2^21 ) )   n = 21   d_n = -1 
assign v[4'b0011] [22] = 22'h 000000;  // -0.0000000000000000 = 2^(22+1) *  0 * atan( 1 / ( -1 + 2^22 ) )   n = 22   d_n = -1 
assign v[4'b0011] [23] = 22'h 000000;  // -0.0000000000000000 = 2^(23+1) *  0 * atan( 1 / ( -1 + 2^23 ) )   n = 23   d_n = -1 
assign v[4'b0011] [24] = 22'h 000000;  // -0.0000000000000000 = 2^(24+1) *  0 * atan( 1 / ( -1 + 2^24 ) )   n = 24   d_n = -1 
assign v[4'b0011] [25] = 22'h 000000;  // -0.0000000000000000 = 2^(25+1) *  0 * atan( 1 / ( -1 + 2^25 ) )   n = 25   d_n = -1 
assign v[4'b0011] [26] = 22'h 000000;  // -0.0000000000000000 = 2^(26+1) *  0 * atan( 1 / ( -1 + 2^26 ) )   n = 26   d_n = -1 
assign v[4'b0011] [27] = 22'h 000000;  // -0.0000000000000000 = 2^(27+1) *  0 * atan( 1 / ( -1 + 2^27 ) )   n = 27   d_n = -1 
assign v[4'b0011] [28] = 22'h 000000;  // -0.0000000000000000 = 2^(28+1) *  0 * atan( 1 / ( -1 + 2^28 ) )   n = 28   d_n = -1 
assign v[4'b0011] [29] = 22'h 000000;  // -0.0000000000000000 = 2^(29+1) *  0 * atan( 1 / ( -1 + 2^29 ) )   n = 29   d_n = -1 
assign v[4'b0011] [30] = 22'h 000000;  // -0.0000000000000000 = 2^(30+1) *  0 * atan( 1 / ( -1 + 2^30 ) )   n = 30   d_n = -1 
assign v[4'b0011] [31] = 22'h 000000;  // -0.0000000000000000 = 2^(31+1) *  0 * atan( 1 / ( -1 + 2^31 ) )   n = 31   d_n = -1 
assign v[4'b0011] [32] = 22'h 000000;  // -0.0000000000000000 = 2^(32+1) *  0 * atan( 1 / ( -1 + 2^32 ) )   n = 32   d_n = -1 
assign v[4'b0011] [33] = 22'h 000000;  // -0.0000000000000000 = 2^(33+1) *  0 * atan( 1 / ( -1 + 2^33 ) )   n = 33   d_n = -1 
assign v[4'b0011] [34] = 22'h 000000;  // -0.0000000000000000 = 2^(34+1) *  0 * atan( 1 / ( -1 + 2^34 ) )   n = 34   d_n = -1 
assign v[4'b0011] [35] = 22'h 000000;  // -0.0000000000000000 = 2^(35+1) *  0 * atan( 1 / ( -1 + 2^35 ) )   n = 35   d_n = -1 
assign v[4'b0011] [36] = 22'h 000000;  // -0.0000000000000000 = 2^(36+1) *  0 * atan( 1 / ( -1 + 2^36 ) )   n = 36   d_n = -1 
assign v[4'b0011] [37] = 22'h 000000;  // -0.0000000000000000 = 2^(37+1) *  0 * atan( 1 / ( -1 + 2^37 ) )   n = 37   d_n = -1 
assign v[4'b0011] [38] = 22'h 000000;  // -0.0000000000000000 = 2^(38+1) *  0 * atan( 1 / ( -1 + 2^38 ) )   n = 38   d_n = -1 
assign v[4'b0011] [39] = 22'h 000000;  // -0.0000000000000000 = 2^(39+1) *  0 * atan( 1 / ( -1 + 2^39 ) )   n = 39   d_n = -1 
assign v[4'b0011] [40] = 22'h 000000;  // -0.0000000000000000 = 2^(40+1) *  0 * atan( 1 / ( -1 + 2^40 ) )   n = 40   d_n = -1 
assign v[4'b0011] [41] = 22'h 000000;  // -0.0000000000000000 = 2^(41+1) *  0 * atan( 1 / ( -1 + 2^41 ) )   n = 41   d_n = -1 
assign v[4'b0011] [42] = 22'h 000000;  // -0.0000000000000000 = 2^(42+1) *  0 * atan( 1 / ( -1 + 2^42 ) )   n = 42   d_n = -1 
assign v[4'b0011] [43] = 22'h 000000;  // -0.0000000000000000 = 2^(43+1) *  0 * atan( 1 / ( -1 + 2^43 ) )   n = 43   d_n = -1 
assign v[4'b0011] [44] = 22'h 000000;  // -0.0000000000000000 = 2^(44+1) *  0 * atan( 1 / ( -1 + 2^44 ) )   n = 44   d_n = -1 
assign v[4'b0011] [45] = 22'h 000000;  // -0.0000000000000000 = 2^(45+1) *  0 * atan( 1 / ( -1 + 2^45 ) )   n = 45   d_n = -1 
assign v[4'b0011] [46] = 22'h 000000;  // -0.0000000000000000 = 2^(46+1) *  0 * atan( 1 / ( -1 + 2^46 ) )   n = 46   d_n = -1 
assign v[4'b0011] [47] = 22'h 000000;  // -0.0000000000000000 = 2^(47+1) *  0 * atan( 1 / ( -1 + 2^47 ) )   n = 47   d_n = -1 
assign v[4'b0011] [48] = 22'h 000000;  // -0.0000000000000000 = 2^(48+1) *  0 * atan( 1 / ( -1 + 2^48 ) )   n = 48   d_n = -1 
assign v[4'b0011] [49] = 22'h 000000;  // -0.0000000000000000 = 2^(49+1) *  0 * atan( 1 / ( -1 + 2^49 ) )   n = 49   d_n = -1 
assign v[4'b0011] [50] = 22'h 000000;  // -0.0000000000000000 = 2^(50+1) *  0 * atan( 1 / ( -1 + 2^50 ) )   n = 50   d_n = -1 
assign v[4'b0011] [51] = 22'h 000000;  // -0.0000000000000000 = 2^(51+1) *  0 * atan( 1 / ( -1 + 2^51 ) )   n = 51   d_n = -1 
assign v[4'b0011] [52] = 22'h 000000;  // -0.0000000000000000 = 2^(52+1) *  0 * atan( 1 / ( -1 + 2^52 ) )   n = 52   d_n = -1 
assign v[4'b0011] [53] = 22'h 000000;  // -0.0000000000000000 = 2^(53+1) *  0 * atan( 1 / ( -1 + 2^53 ) )   n = 53   d_n = -1 
assign v[4'b0011] [54] = 22'h 000000;  // -0.0000000000000000 = 2^(54+1) *  0 * atan( 1 / ( -1 + 2^54 ) )   n = 54   d_n = -1 
assign v[4'b0011] [55] = 22'h 000000;  // -0.0000000000000000 = 2^(55+1) *  0 * atan( 1 / ( -1 + 2^55 ) )   n = 55   d_n = -1 
assign v[4'b0011] [56] = 22'h 000000;  // -0.0000000000000000 = 2^(56+1) *  0 * atan( 1 / ( -1 + 2^56 ) )   n = 56   d_n = -1 
assign v[4'b0011] [57] = 22'h 000000;  // -0.0000000000000000 = 2^(57+1) *  0 * atan( 1 / ( -1 + 2^57 ) )   n = 57   d_n = -1 
assign v[4'b0011] [58] = 22'h 000000;  // -0.0000000000000000 = 2^(58+1) *  0 * atan( 1 / ( -1 + 2^58 ) )   n = 58   d_n = -1 
assign v[4'b0011] [59] = 22'h 000000;  // -0.0000000000000000 = 2^(59+1) *  0 * atan( 1 / ( -1 + 2^59 ) )   n = 59   d_n = -1 
assign v[4'b0011] [60] = 22'h 000000;  // -0.0000000000000000 = 2^(60+1) *  0 * atan( 1 / ( -1 + 2^60 ) )   n = 60   d_n = -1 
assign v[4'b0011] [61] = 22'h 000000;  // -0.0000000000000000 = 2^(61+1) *  0 * atan( 1 / ( -1 + 2^61 ) )   n = 61   d_n = -1 
assign v[4'b0011] [62] = 22'h 000000;  // -0.0000000000000000 = 2^(62+1) *  0 * atan( 1 / ( -1 + 2^62 ) )   n = 62   d_n = -1 
assign v[4'b0011] [63] = 22'h 000000;  // -0.0000000000000000 = 2^(63+1) *  0 * atan( 1 / ( -1 + 2^63 ) )   n = 63   d_n = -1 
assign v[4'b0011] [64] = 22'h 000000;  // -0.0000000000000000 = 2^(64+1) *  0 * atan( 1 / ( -1 + 2^64 ) )   n = 64   d_n = -1 
assign v[4'b0100] [01] = 22'h 0001DA;  // +1.8545904360032244 = 2^(1+1) *  1 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = 0+1i 
assign v[4'b0100] [02] = 22'h 0001F5;  // +1.9598293050149131 = 2^(2+1) *  1 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = 0+1i 
assign v[4'b0100] [03] = 22'h 0001FD;  // +1.9896799127481830 = 2^(3+1) *  1 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = 0+1i 
assign v[4'b0100] [04] = 22'h 0001FF;  // +1.9974019198706352 = 2^(4+1) *  1 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = 0+1i 
assign v[4'b0100] [05] = 22'h 0001FF;  // +1.9993493395371698 = 2^(5+1) *  1 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = 0+1i 
assign v[4'b0100] [06] = 22'h 0001FF;  // +1.9998372634210344 = 2^(6+1) *  1 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = 0+1i 
assign v[4'b0100] [07] = 22'h 0001FF;  // +1.9999593113858845 = 2^(7+1) *  1 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = 0+1i 
assign v[4'b0100] [08] = 22'h 0001FF;  // +1.9999898275670895 = 2^(8+1) *  1 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = 0+1i 
assign v[4'b0100] [09] = 22'h 0001FF;  // +1.9999974568743104 = 2^(9+1) *  1 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = 0+1i 
assign v[4'b0100] [10] = 22'h 0001FF;  // +1.9999993642174863 = 2^(10+1) *  1 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = 0+1i 
assign v[4'b0100] [11] = 22'h 0001FF;  // +1.9999998410543034 = 2^(11+1) *  1 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = 0+1i 
assign v[4'b0100] [12] = 22'h 0001FF;  // +1.9999999602635716 = 2^(12+1) *  1 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = 0+1i 
assign v[4'b0100] [13] = 22'h 0001FF;  // +1.9999999900658927 = 2^(13+1) *  1 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = 0+1i 
assign v[4'b0100] [14] = 22'h 0001FF;  // +1.9999999975164731 = 2^(14+1) *  1 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = 0+1i 
assign v[4'b0100] [15] = 22'h 0001FF;  // +1.9999999993791182 = 2^(15+1) *  1 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = 0+1i 
assign v[4'b0100] [16] = 22'h 0001FF;  // +1.9999999998447795 = 2^(16+1) *  1 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = 0+1i 
assign v[4'b0100] [17] = 22'h 0001FF;  // +1.9999999999611948 = 2^(17+1) *  1 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = 0+1i 
assign v[4'b0100] [18] = 22'h 0001FF;  // +1.9999999999902986 = 2^(18+1) *  1 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = 0+1i 
assign v[4'b0100] [19] = 22'h 0001FF;  // +1.9999999999975746 = 2^(19+1) *  1 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = 0+1i 
assign v[4'b0100] [20] = 22'h 0001FF;  // +1.9999999999993936 = 2^(20+1) *  1 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = 0+1i 
assign v[4'b0100] [21] = 22'h 0001FF;  // +1.9999999999998483 = 2^(21+1) *  1 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = 0+1i 
assign v[4'b0100] [22] = 22'h 0001FF;  // +1.9999999999999620 = 2^(22+1) *  1 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = 0+1i 
assign v[4'b0100] [23] = 22'h 0001FF;  // +1.9999999999999905 = 2^(23+1) *  1 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = 0+1i 
assign v[4'b0100] [24] = 22'h 0001FF;  // +1.9999999999999976 = 2^(24+1) *  1 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = 0+1i 
assign v[4'b0100] [25] = 22'h 0001FF;  // +1.9999999999999993 = 2^(25+1) *  1 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = 0+1i 
assign v[4'b0100] [26] = 22'h 0001FF;  // +1.9999999999999998 = 2^(26+1) *  1 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = 0+1i 
assign v[4'b0100] [27] = 22'h 000200;  // +2.0000000000000000 = 2^(27+1) *  1 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = 0+1i 
assign v[4'b0100] [28] = 22'h 000200;  // +2.0000000000000000 = 2^(28+1) *  1 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = 0+1i 
assign v[4'b0100] [29] = 22'h 000200;  // +2.0000000000000000 = 2^(29+1) *  1 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = 0+1i 
assign v[4'b0100] [30] = 22'h 000200;  // +2.0000000000000000 = 2^(30+1) *  1 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = 0+1i 
assign v[4'b0100] [31] = 22'h 000200;  // +2.0000000000000000 = 2^(31+1) *  1 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = 0+1i 
assign v[4'b0100] [32] = 22'h 000200;  // +2.0000000000000000 = 2^(32+1) *  1 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = 0+1i 
assign v[4'b0100] [33] = 22'h 000200;  // +2.0000000000000000 = 2^(33+1) *  1 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = 0+1i 
assign v[4'b0100] [34] = 22'h 000200;  // +2.0000000000000000 = 2^(34+1) *  1 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = 0+1i 
assign v[4'b0100] [35] = 22'h 000200;  // +2.0000000000000000 = 2^(35+1) *  1 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = 0+1i 
assign v[4'b0100] [36] = 22'h 000200;  // +2.0000000000000000 = 2^(36+1) *  1 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = 0+1i 
assign v[4'b0100] [37] = 22'h 000200;  // +2.0000000000000000 = 2^(37+1) *  1 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = 0+1i 
assign v[4'b0100] [38] = 22'h 000200;  // +2.0000000000000000 = 2^(38+1) *  1 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = 0+1i 
assign v[4'b0100] [39] = 22'h 000200;  // +2.0000000000000000 = 2^(39+1) *  1 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = 0+1i 
assign v[4'b0100] [40] = 22'h 000200;  // +2.0000000000000000 = 2^(40+1) *  1 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = 0+1i 
assign v[4'b0100] [41] = 22'h 000200;  // +2.0000000000000000 = 2^(41+1) *  1 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = 0+1i 
assign v[4'b0100] [42] = 22'h 000200;  // +2.0000000000000000 = 2^(42+1) *  1 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = 0+1i 
assign v[4'b0100] [43] = 22'h 000200;  // +2.0000000000000000 = 2^(43+1) *  1 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = 0+1i 
assign v[4'b0100] [44] = 22'h 000200;  // +2.0000000000000000 = 2^(44+1) *  1 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = 0+1i 
assign v[4'b0100] [45] = 22'h 000200;  // +2.0000000000000000 = 2^(45+1) *  1 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = 0+1i 
assign v[4'b0100] [46] = 22'h 000200;  // +2.0000000000000000 = 2^(46+1) *  1 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = 0+1i 
assign v[4'b0100] [47] = 22'h 000200;  // +2.0000000000000000 = 2^(47+1) *  1 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = 0+1i 
assign v[4'b0100] [48] = 22'h 000200;  // +2.0000000000000000 = 2^(48+1) *  1 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = 0+1i 
assign v[4'b0100] [49] = 22'h 000200;  // +2.0000000000000000 = 2^(49+1) *  1 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = 0+1i 
assign v[4'b0100] [50] = 22'h 000200;  // +2.0000000000000000 = 2^(50+1) *  1 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = 0+1i 
assign v[4'b0100] [51] = 22'h 000200;  // +2.0000000000000000 = 2^(51+1) *  1 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = 0+1i 
assign v[4'b0100] [52] = 22'h 000200;  // +2.0000000000000000 = 2^(52+1) *  1 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = 0+1i 
assign v[4'b0100] [53] = 22'h 000200;  // +2.0000000000000000 = 2^(53+1) *  1 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = 0+1i 
assign v[4'b0100] [54] = 22'h 000200;  // +2.0000000000000000 = 2^(54+1) *  1 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = 0+1i 
assign v[4'b0100] [55] = 22'h 000200;  // +2.0000000000000000 = 2^(55+1) *  1 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = 0+1i 
assign v[4'b0100] [56] = 22'h 000200;  // +2.0000000000000000 = 2^(56+1) *  1 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = 0+1i 
assign v[4'b0100] [57] = 22'h 000200;  // +2.0000000000000000 = 2^(57+1) *  1 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = 0+1i 
assign v[4'b0100] [58] = 22'h 000200;  // +2.0000000000000000 = 2^(58+1) *  1 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = 0+1i 
assign v[4'b0100] [59] = 22'h 000200;  // +2.0000000000000000 = 2^(59+1) *  1 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = 0+1i 
assign v[4'b0100] [60] = 22'h 000200;  // +2.0000000000000000 = 2^(60+1) *  1 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = 0+1i 
assign v[4'b0100] [61] = 22'h 000200;  // +2.0000000000000000 = 2^(61+1) *  1 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = 0+1i 
assign v[4'b0100] [62] = 22'h 000200;  // +2.0000000000000000 = 2^(62+1) *  1 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = 0+1i 
assign v[4'b0100] [63] = 22'h 000200;  // +2.0000000000000000 = 2^(63+1) *  1 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = 0+1i 
assign v[4'b0100] [64] = 22'h 000200;  // +2.0000000000000000 = 2^(64+1) *  1 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = 0+1i 
assign v[4'b0101] [01] = 22'h 000149;  // +1.2870022175865687 = 2^(1+1) *  1 * atan( 1 / (  1 + 2^1 ) )   n =  1   d_n = 1+1i 
assign v[4'b0101] [02] = 22'h 000194;  // +1.5791644787990460 = 2^(2+1) *  1 * atan( 1 / (  1 + 2^2 ) )   n =  2   d_n = 1+1i 
assign v[4'b0101] [03] = 22'h 0001C5;  // +1.7705155387823304 = 2^(3+1) *  1 * atan( 1 / (  1 + 2^3 ) )   n =  3   d_n = 1+1i 
assign v[4'b0101] [04] = 22'h 0001E1;  // +1.8801863269031263 = 2^(4+1) *  1 * atan( 1 / (  1 + 2^4 ) )   n =  4   d_n = 1+1i 
assign v[4'b0101] [05] = 22'h 0001F0;  // +1.9388006348016065 = 2^(5+1) *  1 * atan( 1 / (  1 + 2^5 ) )   n =  5   d_n = 1+1i 
assign v[4'b0101] [06] = 22'h 0001F8;  // +1.9690754279161793 = 2^(6+1) *  1 * atan( 1 / (  1 + 2^6 ) )   n =  6   d_n = 1+1i 
assign v[4'b0101] [07] = 22'h 0001FC;  // +1.9844563743249595 = 2^(7+1) *  1 * atan( 1 / (  1 + 2^7 ) )   n =  7   d_n = 1+1i 
assign v[4'b0101] [08] = 22'h 0001FE;  // +1.9922078446819715 = 2^(8+1) *  1 * atan( 1 / (  1 + 2^8 ) )   n =  8   d_n = 1+1i 
assign v[4'b0101] [09] = 22'h 0001FF;  // +1.9960988362398133 = 2^(9+1) *  1 * atan( 1 / (  1 + 2^9 ) )   n =  9   d_n = 1+1i 
assign v[4'b0101] [10] = 22'h 0001FF;  // +1.9980481465643023 = 2^(10+1) *  1 * atan( 1 / (  1 + 2^10 ) )   n = 10   d_n = 1+1i 
assign v[4'b0101] [11] = 22'h 0001FF;  // +1.9990237553913479 = 2^(11+1) *  1 * atan( 1 / (  1 + 2^11 ) )   n = 11   d_n = 1+1i 
assign v[4'b0101] [12] = 22'h 0001FF;  // +1.9995117982228541 = 2^(12+1) *  1 * atan( 1 / (  1 + 2^12 ) )   n = 12   d_n = 1+1i 
assign v[4'b0101] [13] = 22'h 0001FF;  // +1.9997558792432146 = 2^(13+1) *  1 * atan( 1 / (  1 + 2^13 ) )   n = 13   d_n = 1+1i 
assign v[4'b0101] [14] = 22'h 0001FF;  // +1.9998779346545537 = 2^(14+1) *  1 * atan( 1 / (  1 + 2^14 ) )   n = 14   d_n = 1+1i 
assign v[4'b0101] [15] = 22'h 0001FF;  // +1.9999389660855134 = 2^(15+1) *  1 * atan( 1 / (  1 + 2^15 ) )   n = 15   d_n = 1+1i 
assign v[4'b0101] [16] = 22'h 0001FF;  // +1.9999694827323158 = 2^(16+1) *  1 * atan( 1 / (  1 + 2^16 ) )   n = 16   d_n = 1+1i 
assign v[4'b0101] [17] = 22'h 0001FF;  // +1.9999847412885476 = 2^(17+1) *  1 * atan( 1 / (  1 + 2^17 ) )   n = 17   d_n = 1+1i 
assign v[4'b0101] [18] = 22'h 0001FF;  // +1.9999923706248712 = 2^(18+1) *  1 * atan( 1 / (  1 + 2^18 ) )   n = 18   d_n = 1+1i 
assign v[4'b0101] [19] = 22'h 0001FF;  // +1.9999961853075849 = 2^(19+1) *  1 * atan( 1 / (  1 + 2^19 ) )   n = 19   d_n = 1+1i 
assign v[4'b0101] [20] = 22'h 0001FF;  // +1.9999980926525798 = 2^(20+1) *  1 * atan( 1 / (  1 + 2^20 ) )   n = 20   d_n = 1+1i 
assign v[4'b0101] [21] = 22'h 0001FF;  // +1.9999990463259867 = 2^(21+1) *  1 * atan( 1 / (  1 + 2^21 ) )   n = 21   d_n = 1+1i 
assign v[4'b0101] [22] = 22'h 0001FF;  // +1.9999995231629175 = 2^(22+1) *  1 * atan( 1 / (  1 + 2^22 ) )   n = 22   d_n = 1+1i 
assign v[4'b0101] [23] = 22'h 0001FF;  // +1.9999997615814398 = 2^(23+1) *  1 * atan( 1 / (  1 + 2^23 ) )   n = 23   d_n = 1+1i 
assign v[4'b0101] [24] = 22'h 0001FF;  // +1.9999998807907151 = 2^(24+1) *  1 * atan( 1 / (  1 + 2^24 ) )   n = 24   d_n = 1+1i 
assign v[4'b0101] [25] = 22'h 0001FF;  // +1.9999999403953563 = 2^(25+1) *  1 * atan( 1 / (  1 + 2^25 ) )   n = 25   d_n = 1+1i 
assign v[4'b0101] [26] = 22'h 0001FF;  // +1.9999999701976778 = 2^(26+1) *  1 * atan( 1 / (  1 + 2^26 ) )   n = 26   d_n = 1+1i 
assign v[4'b0101] [27] = 22'h 0001FF;  // +1.9999999850988388 = 2^(27+1) *  1 * atan( 1 / (  1 + 2^27 ) )   n = 27   d_n = 1+1i 
assign v[4'b0101] [28] = 22'h 0001FF;  // +1.9999999925494194 = 2^(28+1) *  1 * atan( 1 / (  1 + 2^28 ) )   n = 28   d_n = 1+1i 
assign v[4'b0101] [29] = 22'h 0001FF;  // +1.9999999962747097 = 2^(29+1) *  1 * atan( 1 / (  1 + 2^29 ) )   n = 29   d_n = 1+1i 
assign v[4'b0101] [30] = 22'h 0001FF;  // +1.9999999981373549 = 2^(30+1) *  1 * atan( 1 / (  1 + 2^30 ) )   n = 30   d_n = 1+1i 
assign v[4'b0101] [31] = 22'h 0001FF;  // +1.9999999990686774 = 2^(31+1) *  1 * atan( 1 / (  1 + 2^31 ) )   n = 31   d_n = 1+1i 
assign v[4'b0101] [32] = 22'h 0001FF;  // +1.9999999995343387 = 2^(32+1) *  1 * atan( 1 / (  1 + 2^32 ) )   n = 32   d_n = 1+1i 
assign v[4'b0101] [33] = 22'h 0001FF;  // +1.9999999997671694 = 2^(33+1) *  1 * atan( 1 / (  1 + 2^33 ) )   n = 33   d_n = 1+1i 
assign v[4'b0101] [34] = 22'h 0001FF;  // +1.9999999998835847 = 2^(34+1) *  1 * atan( 1 / (  1 + 2^34 ) )   n = 34   d_n = 1+1i 
assign v[4'b0101] [35] = 22'h 0001FF;  // +1.9999999999417923 = 2^(35+1) *  1 * atan( 1 / (  1 + 2^35 ) )   n = 35   d_n = 1+1i 
assign v[4'b0101] [36] = 22'h 0001FF;  // +1.9999999999708962 = 2^(36+1) *  1 * atan( 1 / (  1 + 2^36 ) )   n = 36   d_n = 1+1i 
assign v[4'b0101] [37] = 22'h 0001FF;  // +1.9999999999854481 = 2^(37+1) *  1 * atan( 1 / (  1 + 2^37 ) )   n = 37   d_n = 1+1i 
assign v[4'b0101] [38] = 22'h 0001FF;  // +1.9999999999927240 = 2^(38+1) *  1 * atan( 1 / (  1 + 2^38 ) )   n = 38   d_n = 1+1i 
assign v[4'b0101] [39] = 22'h 0001FF;  // +1.9999999999963620 = 2^(39+1) *  1 * atan( 1 / (  1 + 2^39 ) )   n = 39   d_n = 1+1i 
assign v[4'b0101] [40] = 22'h 0001FF;  // +1.9999999999981810 = 2^(40+1) *  1 * atan( 1 / (  1 + 2^40 ) )   n = 40   d_n = 1+1i 
assign v[4'b0101] [41] = 22'h 0001FF;  // +1.9999999999990905 = 2^(41+1) *  1 * atan( 1 / (  1 + 2^41 ) )   n = 41   d_n = 1+1i 
assign v[4'b0101] [42] = 22'h 0001FF;  // +1.9999999999995453 = 2^(42+1) *  1 * atan( 1 / (  1 + 2^42 ) )   n = 42   d_n = 1+1i 
assign v[4'b0101] [43] = 22'h 0001FF;  // +1.9999999999997726 = 2^(43+1) *  1 * atan( 1 / (  1 + 2^43 ) )   n = 43   d_n = 1+1i 
assign v[4'b0101] [44] = 22'h 0001FF;  // +1.9999999999998863 = 2^(44+1) *  1 * atan( 1 / (  1 + 2^44 ) )   n = 44   d_n = 1+1i 
assign v[4'b0101] [45] = 22'h 0001FF;  // +1.9999999999999432 = 2^(45+1) *  1 * atan( 1 / (  1 + 2^45 ) )   n = 45   d_n = 1+1i 
assign v[4'b0101] [46] = 22'h 0001FF;  // +1.9999999999999716 = 2^(46+1) *  1 * atan( 1 / (  1 + 2^46 ) )   n = 46   d_n = 1+1i 
assign v[4'b0101] [47] = 22'h 0001FF;  // +1.9999999999999858 = 2^(47+1) *  1 * atan( 1 / (  1 + 2^47 ) )   n = 47   d_n = 1+1i 
assign v[4'b0101] [48] = 22'h 0001FF;  // +1.9999999999999929 = 2^(48+1) *  1 * atan( 1 / (  1 + 2^48 ) )   n = 48   d_n = 1+1i 
assign v[4'b0101] [49] = 22'h 0001FF;  // +1.9999999999999964 = 2^(49+1) *  1 * atan( 1 / (  1 + 2^49 ) )   n = 49   d_n = 1+1i 
assign v[4'b0101] [50] = 22'h 0001FF;  // +1.9999999999999982 = 2^(50+1) *  1 * atan( 1 / (  1 + 2^50 ) )   n = 50   d_n = 1+1i 
assign v[4'b0101] [51] = 22'h 0001FF;  // +1.9999999999999991 = 2^(51+1) *  1 * atan( 1 / (  1 + 2^51 ) )   n = 51   d_n = 1+1i 
assign v[4'b0101] [52] = 22'h 0001FF;  // +1.9999999999999996 = 2^(52+1) *  1 * atan( 1 / (  1 + 2^52 ) )   n = 52   d_n = 1+1i 
assign v[4'b0101] [53] = 22'h 000200;  // +2.0000000000000000 = 2^(53+1) *  1 * atan( 1 / (  1 + 2^53 ) )   n = 53   d_n = 1+1i 
assign v[4'b0101] [54] = 22'h 000200;  // +2.0000000000000000 = 2^(54+1) *  1 * atan( 1 / (  1 + 2^54 ) )   n = 54   d_n = 1+1i 
assign v[4'b0101] [55] = 22'h 000200;  // +2.0000000000000000 = 2^(55+1) *  1 * atan( 1 / (  1 + 2^55 ) )   n = 55   d_n = 1+1i 
assign v[4'b0101] [56] = 22'h 000200;  // +2.0000000000000000 = 2^(56+1) *  1 * atan( 1 / (  1 + 2^56 ) )   n = 56   d_n = 1+1i 
assign v[4'b0101] [57] = 22'h 000200;  // +2.0000000000000000 = 2^(57+1) *  1 * atan( 1 / (  1 + 2^57 ) )   n = 57   d_n = 1+1i 
assign v[4'b0101] [58] = 22'h 000200;  // +2.0000000000000000 = 2^(58+1) *  1 * atan( 1 / (  1 + 2^58 ) )   n = 58   d_n = 1+1i 
assign v[4'b0101] [59] = 22'h 000200;  // +2.0000000000000000 = 2^(59+1) *  1 * atan( 1 / (  1 + 2^59 ) )   n = 59   d_n = 1+1i 
assign v[4'b0101] [60] = 22'h 000200;  // +2.0000000000000000 = 2^(60+1) *  1 * atan( 1 / (  1 + 2^60 ) )   n = 60   d_n = 1+1i 
assign v[4'b0101] [61] = 22'h 000200;  // +2.0000000000000000 = 2^(61+1) *  1 * atan( 1 / (  1 + 2^61 ) )   n = 61   d_n = 1+1i 
assign v[4'b0101] [62] = 22'h 000200;  // +2.0000000000000000 = 2^(62+1) *  1 * atan( 1 / (  1 + 2^62 ) )   n = 62   d_n = 1+1i 
assign v[4'b0101] [63] = 22'h 000200;  // +2.0000000000000000 = 2^(63+1) *  1 * atan( 1 / (  1 + 2^63 ) )   n = 63   d_n = 1+1i 
assign v[4'b0101] [64] = 22'h 000200;  // +2.0000000000000000 = 2^(64+1) *  1 * atan( 1 / (  1 + 2^64 ) )   n = 64   d_n = 1+1i 
assign v[4'b0110] [01] = 22'h 0001DA;  // +1.8545904360032244 = 2^(1+1) *  1 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = 0+1i 
assign v[4'b0110] [02] = 22'h 0001F5;  // +1.9598293050149131 = 2^(2+1) *  1 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = 0+1i 
assign v[4'b0110] [03] = 22'h 0001FD;  // +1.9896799127481830 = 2^(3+1) *  1 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = 0+1i 
assign v[4'b0110] [04] = 22'h 0001FF;  // +1.9974019198706352 = 2^(4+1) *  1 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = 0+1i 
assign v[4'b0110] [05] = 22'h 0001FF;  // +1.9993493395371698 = 2^(5+1) *  1 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = 0+1i 
assign v[4'b0110] [06] = 22'h 0001FF;  // +1.9998372634210344 = 2^(6+1) *  1 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = 0+1i 
assign v[4'b0110] [07] = 22'h 0001FF;  // +1.9999593113858845 = 2^(7+1) *  1 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = 0+1i 
assign v[4'b0110] [08] = 22'h 0001FF;  // +1.9999898275670895 = 2^(8+1) *  1 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = 0+1i 
assign v[4'b0110] [09] = 22'h 0001FF;  // +1.9999974568743104 = 2^(9+1) *  1 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = 0+1i 
assign v[4'b0110] [10] = 22'h 0001FF;  // +1.9999993642174863 = 2^(10+1) *  1 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = 0+1i 
assign v[4'b0110] [11] = 22'h 0001FF;  // +1.9999998410543034 = 2^(11+1) *  1 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = 0+1i 
assign v[4'b0110] [12] = 22'h 0001FF;  // +1.9999999602635716 = 2^(12+1) *  1 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = 0+1i 
assign v[4'b0110] [13] = 22'h 0001FF;  // +1.9999999900658927 = 2^(13+1) *  1 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = 0+1i 
assign v[4'b0110] [14] = 22'h 0001FF;  // +1.9999999975164731 = 2^(14+1) *  1 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = 0+1i 
assign v[4'b0110] [15] = 22'h 0001FF;  // +1.9999999993791182 = 2^(15+1) *  1 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = 0+1i 
assign v[4'b0110] [16] = 22'h 0001FF;  // +1.9999999998447795 = 2^(16+1) *  1 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = 0+1i 
assign v[4'b0110] [17] = 22'h 0001FF;  // +1.9999999999611948 = 2^(17+1) *  1 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = 0+1i 
assign v[4'b0110] [18] = 22'h 0001FF;  // +1.9999999999902986 = 2^(18+1) *  1 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = 0+1i 
assign v[4'b0110] [19] = 22'h 0001FF;  // +1.9999999999975746 = 2^(19+1) *  1 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = 0+1i 
assign v[4'b0110] [20] = 22'h 0001FF;  // +1.9999999999993936 = 2^(20+1) *  1 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = 0+1i 
assign v[4'b0110] [21] = 22'h 0001FF;  // +1.9999999999998483 = 2^(21+1) *  1 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = 0+1i 
assign v[4'b0110] [22] = 22'h 0001FF;  // +1.9999999999999620 = 2^(22+1) *  1 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = 0+1i 
assign v[4'b0110] [23] = 22'h 0001FF;  // +1.9999999999999905 = 2^(23+1) *  1 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = 0+1i 
assign v[4'b0110] [24] = 22'h 0001FF;  // +1.9999999999999976 = 2^(24+1) *  1 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = 0+1i 
assign v[4'b0110] [25] = 22'h 0001FF;  // +1.9999999999999993 = 2^(25+1) *  1 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = 0+1i 
assign v[4'b0110] [26] = 22'h 0001FF;  // +1.9999999999999998 = 2^(26+1) *  1 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = 0+1i 
assign v[4'b0110] [27] = 22'h 000200;  // +2.0000000000000000 = 2^(27+1) *  1 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = 0+1i 
assign v[4'b0110] [28] = 22'h 000200;  // +2.0000000000000000 = 2^(28+1) *  1 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = 0+1i 
assign v[4'b0110] [29] = 22'h 000200;  // +2.0000000000000000 = 2^(29+1) *  1 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = 0+1i 
assign v[4'b0110] [30] = 22'h 000200;  // +2.0000000000000000 = 2^(30+1) *  1 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = 0+1i 
assign v[4'b0110] [31] = 22'h 000200;  // +2.0000000000000000 = 2^(31+1) *  1 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = 0+1i 
assign v[4'b0110] [32] = 22'h 000200;  // +2.0000000000000000 = 2^(32+1) *  1 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = 0+1i 
assign v[4'b0110] [33] = 22'h 000200;  // +2.0000000000000000 = 2^(33+1) *  1 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = 0+1i 
assign v[4'b0110] [34] = 22'h 000200;  // +2.0000000000000000 = 2^(34+1) *  1 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = 0+1i 
assign v[4'b0110] [35] = 22'h 000200;  // +2.0000000000000000 = 2^(35+1) *  1 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = 0+1i 
assign v[4'b0110] [36] = 22'h 000200;  // +2.0000000000000000 = 2^(36+1) *  1 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = 0+1i 
assign v[4'b0110] [37] = 22'h 000200;  // +2.0000000000000000 = 2^(37+1) *  1 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = 0+1i 
assign v[4'b0110] [38] = 22'h 000200;  // +2.0000000000000000 = 2^(38+1) *  1 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = 0+1i 
assign v[4'b0110] [39] = 22'h 000200;  // +2.0000000000000000 = 2^(39+1) *  1 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = 0+1i 
assign v[4'b0110] [40] = 22'h 000200;  // +2.0000000000000000 = 2^(40+1) *  1 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = 0+1i 
assign v[4'b0110] [41] = 22'h 000200;  // +2.0000000000000000 = 2^(41+1) *  1 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = 0+1i 
assign v[4'b0110] [42] = 22'h 000200;  // +2.0000000000000000 = 2^(42+1) *  1 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = 0+1i 
assign v[4'b0110] [43] = 22'h 000200;  // +2.0000000000000000 = 2^(43+1) *  1 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = 0+1i 
assign v[4'b0110] [44] = 22'h 000200;  // +2.0000000000000000 = 2^(44+1) *  1 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = 0+1i 
assign v[4'b0110] [45] = 22'h 000200;  // +2.0000000000000000 = 2^(45+1) *  1 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = 0+1i 
assign v[4'b0110] [46] = 22'h 000200;  // +2.0000000000000000 = 2^(46+1) *  1 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = 0+1i 
assign v[4'b0110] [47] = 22'h 000200;  // +2.0000000000000000 = 2^(47+1) *  1 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = 0+1i 
assign v[4'b0110] [48] = 22'h 000200;  // +2.0000000000000000 = 2^(48+1) *  1 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = 0+1i 
assign v[4'b0110] [49] = 22'h 000200;  // +2.0000000000000000 = 2^(49+1) *  1 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = 0+1i 
assign v[4'b0110] [50] = 22'h 000200;  // +2.0000000000000000 = 2^(50+1) *  1 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = 0+1i 
assign v[4'b0110] [51] = 22'h 000200;  // +2.0000000000000000 = 2^(51+1) *  1 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = 0+1i 
assign v[4'b0110] [52] = 22'h 000200;  // +2.0000000000000000 = 2^(52+1) *  1 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = 0+1i 
assign v[4'b0110] [53] = 22'h 000200;  // +2.0000000000000000 = 2^(53+1) *  1 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = 0+1i 
assign v[4'b0110] [54] = 22'h 000200;  // +2.0000000000000000 = 2^(54+1) *  1 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = 0+1i 
assign v[4'b0110] [55] = 22'h 000200;  // +2.0000000000000000 = 2^(55+1) *  1 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = 0+1i 
assign v[4'b0110] [56] = 22'h 000200;  // +2.0000000000000000 = 2^(56+1) *  1 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = 0+1i 
assign v[4'b0110] [57] = 22'h 000200;  // +2.0000000000000000 = 2^(57+1) *  1 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = 0+1i 
assign v[4'b0110] [58] = 22'h 000200;  // +2.0000000000000000 = 2^(58+1) *  1 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = 0+1i 
assign v[4'b0110] [59] = 22'h 000200;  // +2.0000000000000000 = 2^(59+1) *  1 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = 0+1i 
assign v[4'b0110] [60] = 22'h 000200;  // +2.0000000000000000 = 2^(60+1) *  1 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = 0+1i 
assign v[4'b0110] [61] = 22'h 000200;  // +2.0000000000000000 = 2^(61+1) *  1 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = 0+1i 
assign v[4'b0110] [62] = 22'h 000200;  // +2.0000000000000000 = 2^(62+1) *  1 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = 0+1i 
assign v[4'b0110] [63] = 22'h 000200;  // +2.0000000000000000 = 2^(63+1) *  1 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = 0+1i 
assign v[4'b0110] [64] = 22'h 000200;  // +2.0000000000000000 = 2^(64+1) *  1 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = 0+1i 
assign v[4'b0111] [01] = 22'h 000324;  // +3.1415926535897931 = 2^(1+1) *  1 * atan( 1 / ( -1 + 2^1 ) )   n =  1   d_n = -1+1i 
assign v[4'b0111] [02] = 22'h 000292;  // +2.5740044351731375 = 2^(2+1) *  1 * atan( 1 / ( -1 + 2^2 ) )   n =  2   d_n = -1+1i 
assign v[4'b0111] [03] = 22'h 000245;  // +2.2703528736666230 = 2^(3+1) *  1 * atan( 1 / ( -1 + 2^3 ) )   n =  3   d_n = -1+1i 
assign v[4'b0111] [04] = 22'h 000221;  // +2.1301812408263618 = 2^(4+1) *  1 * atan( 1 / ( -1 + 2^4 ) )   n =  4   d_n = -1+1i 
assign v[4'b0111] [05] = 22'h 000210;  // +2.0638004758562509 = 2^(5+1) *  1 * atan( 1 / ( -1 + 2^5 ) )   n =  5   d_n = -1+1i 
assign v[4'b0111] [06] = 22'h 000208;  // +2.0315754229491265 = 2^(6+1) *  1 * atan( 1 / ( -1 + 2^6 ) )   n =  6   d_n = -1+1i 
assign v[4'b0111] [07] = 22'h 000204;  // +2.0157063741697390 = 2^(7+1) *  1 * atan( 1 / ( -1 + 2^7 ) )   n =  7   d_n = -1+1i 
assign v[4'b0111] [08] = 22'h 000202;  // +2.0078328446771208 = 2^(8+1) *  1 * atan( 1 / ( -1 + 2^8 ) )   n =  8   d_n = -1+1i 
assign v[4'b0111] [09] = 22'h 000201;  // +2.0039113362396619 = 2^(9+1) *  1 * atan( 1 / ( -1 + 2^9 ) )   n =  9   d_n = -1+1i 
assign v[4'b0111] [10] = 22'h 000200;  // +2.0019543965642979 = 2^(10+1) *  1 * atan( 1 / ( -1 + 2^10 ) )   n = 10   d_n = -1+1i 
assign v[4'b0111] [11] = 22'h 000200;  // +2.0009768803913479 = 2^(11+1) *  1 * atan( 1 / ( -1 + 2^11 ) )   n = 11   d_n = -1+1i 
assign v[4'b0111] [12] = 22'h 000200;  // +2.0004883607228541 = 2^(12+1) *  1 * atan( 1 / ( -1 + 2^12 ) )   n = 12   d_n = -1+1i 
assign v[4'b0111] [13] = 22'h 000200;  // +2.0002441604932146 = 2^(13+1) *  1 * atan( 1 / ( -1 + 2^13 ) )   n = 13   d_n = -1+1i 
assign v[4'b0111] [14] = 22'h 000200;  // +2.0001220752795539 = 2^(14+1) *  1 * atan( 1 / ( -1 + 2^14 ) )   n = 14   d_n = -1+1i 
assign v[4'b0111] [15] = 22'h 000200;  // +2.0000610363980136 = 2^(15+1) *  1 * atan( 1 / ( -1 + 2^15 ) )   n = 15   d_n = -1+1i 
assign v[4'b0111] [16] = 22'h 000200;  // +2.0000305178885660 = 2^(16+1) *  1 * atan( 1 / ( -1 + 2^16 ) )   n = 16   d_n = -1+1i 
assign v[4'b0111] [17] = 22'h 000200;  // +2.0000152588666729 = 2^(17+1) *  1 * atan( 1 / ( -1 + 2^17 ) )   n = 17   d_n = -1+1i 
assign v[4'b0111] [18] = 22'h 000200;  // +2.0000076294139340 = 2^(18+1) *  1 * atan( 1 / ( -1 + 2^18 ) )   n = 18   d_n = -1+1i 
assign v[4'b0111] [19] = 22'h 000200;  // +2.0000038147021164 = 2^(19+1) *  1 * atan( 1 / ( -1 + 2^19 ) )   n = 19   d_n = -1+1i 
assign v[4'b0111] [20] = 22'h 000200;  // +2.0000019073498456 = 2^(20+1) *  1 * atan( 1 / ( -1 + 2^20 ) )   n = 20   d_n = -1+1i 
assign v[4'b0111] [21] = 22'h 000200;  // +2.0000009536746197 = 2^(21+1) *  1 * atan( 1 / ( -1 + 2^21 ) )   n = 21   d_n = -1+1i 
assign v[4'b0111] [22] = 22'h 000200;  // +2.0000004768372341 = 2^(22+1) *  1 * atan( 1 / ( -1 + 2^22 ) )   n = 22   d_n = -1+1i 
assign v[4'b0111] [23] = 22'h 000200;  // +2.0000002384185982 = 2^(23+1) *  1 * atan( 1 / ( -1 + 2^23 ) )   n = 23   d_n = -1+1i 
assign v[4'b0111] [24] = 22'h 000200;  // +2.0000001192092944 = 2^(24+1) *  1 * atan( 1 / ( -1 + 2^24 ) )   n = 24   d_n = -1+1i 
assign v[4'b0111] [25] = 22'h 000200;  // +2.0000000596046461 = 2^(25+1) *  1 * atan( 1 / ( -1 + 2^25 ) )   n = 25   d_n = -1+1i 
assign v[4'b0111] [26] = 22'h 000200;  // +2.0000000298023228 = 2^(26+1) *  1 * atan( 1 / ( -1 + 2^26 ) )   n = 26   d_n = -1+1i 
assign v[4'b0111] [27] = 22'h 000200;  // +2.0000000149011612 = 2^(27+1) *  1 * atan( 1 / ( -1 + 2^27 ) )   n = 27   d_n = -1+1i 
assign v[4'b0111] [28] = 22'h 000200;  // +2.0000000074505806 = 2^(28+1) *  1 * atan( 1 / ( -1 + 2^28 ) )   n = 28   d_n = -1+1i 
assign v[4'b0111] [29] = 22'h 000200;  // +2.0000000037252903 = 2^(29+1) *  1 * atan( 1 / ( -1 + 2^29 ) )   n = 29   d_n = -1+1i 
assign v[4'b0111] [30] = 22'h 000200;  // +2.0000000018626451 = 2^(30+1) *  1 * atan( 1 / ( -1 + 2^30 ) )   n = 30   d_n = -1+1i 
assign v[4'b0111] [31] = 22'h 000200;  // +2.0000000009313226 = 2^(31+1) *  1 * atan( 1 / ( -1 + 2^31 ) )   n = 31   d_n = -1+1i 
assign v[4'b0111] [32] = 22'h 000200;  // +2.0000000004656613 = 2^(32+1) *  1 * atan( 1 / ( -1 + 2^32 ) )   n = 32   d_n = -1+1i 
assign v[4'b0111] [33] = 22'h 000200;  // +2.0000000002328306 = 2^(33+1) *  1 * atan( 1 / ( -1 + 2^33 ) )   n = 33   d_n = -1+1i 
assign v[4'b0111] [34] = 22'h 000200;  // +2.0000000001164153 = 2^(34+1) *  1 * atan( 1 / ( -1 + 2^34 ) )   n = 34   d_n = -1+1i 
assign v[4'b0111] [35] = 22'h 000200;  // +2.0000000000582077 = 2^(35+1) *  1 * atan( 1 / ( -1 + 2^35 ) )   n = 35   d_n = -1+1i 
assign v[4'b0111] [36] = 22'h 000200;  // +2.0000000000291038 = 2^(36+1) *  1 * atan( 1 / ( -1 + 2^36 ) )   n = 36   d_n = -1+1i 
assign v[4'b0111] [37] = 22'h 000200;  // +2.0000000000145519 = 2^(37+1) *  1 * atan( 1 / ( -1 + 2^37 ) )   n = 37   d_n = -1+1i 
assign v[4'b0111] [38] = 22'h 000200;  // +2.0000000000072760 = 2^(38+1) *  1 * atan( 1 / ( -1 + 2^38 ) )   n = 38   d_n = -1+1i 
assign v[4'b0111] [39] = 22'h 000200;  // +2.0000000000036380 = 2^(39+1) *  1 * atan( 1 / ( -1 + 2^39 ) )   n = 39   d_n = -1+1i 
assign v[4'b0111] [40] = 22'h 000200;  // +2.0000000000018190 = 2^(40+1) *  1 * atan( 1 / ( -1 + 2^40 ) )   n = 40   d_n = -1+1i 
assign v[4'b0111] [41] = 22'h 000200;  // +2.0000000000009095 = 2^(41+1) *  1 * atan( 1 / ( -1 + 2^41 ) )   n = 41   d_n = -1+1i 
assign v[4'b0111] [42] = 22'h 000200;  // +2.0000000000004547 = 2^(42+1) *  1 * atan( 1 / ( -1 + 2^42 ) )   n = 42   d_n = -1+1i 
assign v[4'b0111] [43] = 22'h 000200;  // +2.0000000000002274 = 2^(43+1) *  1 * atan( 1 / ( -1 + 2^43 ) )   n = 43   d_n = -1+1i 
assign v[4'b0111] [44] = 22'h 000200;  // +2.0000000000001137 = 2^(44+1) *  1 * atan( 1 / ( -1 + 2^44 ) )   n = 44   d_n = -1+1i 
assign v[4'b0111] [45] = 22'h 000200;  // +2.0000000000000568 = 2^(45+1) *  1 * atan( 1 / ( -1 + 2^45 ) )   n = 45   d_n = -1+1i 
assign v[4'b0111] [46] = 22'h 000200;  // +2.0000000000000284 = 2^(46+1) *  1 * atan( 1 / ( -1 + 2^46 ) )   n = 46   d_n = -1+1i 
assign v[4'b0111] [47] = 22'h 000200;  // +2.0000000000000142 = 2^(47+1) *  1 * atan( 1 / ( -1 + 2^47 ) )   n = 47   d_n = -1+1i 
assign v[4'b0111] [48] = 22'h 000200;  // +2.0000000000000071 = 2^(48+1) *  1 * atan( 1 / ( -1 + 2^48 ) )   n = 48   d_n = -1+1i 
assign v[4'b0111] [49] = 22'h 000200;  // +2.0000000000000036 = 2^(49+1) *  1 * atan( 1 / ( -1 + 2^49 ) )   n = 49   d_n = -1+1i 
assign v[4'b0111] [50] = 22'h 000200;  // +2.0000000000000018 = 2^(50+1) *  1 * atan( 1 / ( -1 + 2^50 ) )   n = 50   d_n = -1+1i 
assign v[4'b0111] [51] = 22'h 000200;  // +2.0000000000000009 = 2^(51+1) *  1 * atan( 1 / ( -1 + 2^51 ) )   n = 51   d_n = -1+1i 
assign v[4'b0111] [52] = 22'h 000200;  // +2.0000000000000004 = 2^(52+1) *  1 * atan( 1 / ( -1 + 2^52 ) )   n = 52   d_n = -1+1i 
assign v[4'b0111] [53] = 22'h 000200;  // +2.0000000000000004 = 2^(53+1) *  1 * atan( 1 / ( -1 + 2^53 ) )   n = 53   d_n = -1+1i 
assign v[4'b0111] [54] = 22'h 000200;  // +2.0000000000000000 = 2^(54+1) *  1 * atan( 1 / ( -1 + 2^54 ) )   n = 54   d_n = -1+1i 
assign v[4'b0111] [55] = 22'h 000200;  // +2.0000000000000000 = 2^(55+1) *  1 * atan( 1 / ( -1 + 2^55 ) )   n = 55   d_n = -1+1i 
assign v[4'b0111] [56] = 22'h 000200;  // +2.0000000000000000 = 2^(56+1) *  1 * atan( 1 / ( -1 + 2^56 ) )   n = 56   d_n = -1+1i 
assign v[4'b0111] [57] = 22'h 000200;  // +2.0000000000000000 = 2^(57+1) *  1 * atan( 1 / ( -1 + 2^57 ) )   n = 57   d_n = -1+1i 
assign v[4'b0111] [58] = 22'h 000200;  // +2.0000000000000000 = 2^(58+1) *  1 * atan( 1 / ( -1 + 2^58 ) )   n = 58   d_n = -1+1i 
assign v[4'b0111] [59] = 22'h 000200;  // +2.0000000000000000 = 2^(59+1) *  1 * atan( 1 / ( -1 + 2^59 ) )   n = 59   d_n = -1+1i 
assign v[4'b0111] [60] = 22'h 000200;  // +2.0000000000000000 = 2^(60+1) *  1 * atan( 1 / ( -1 + 2^60 ) )   n = 60   d_n = -1+1i 
assign v[4'b0111] [61] = 22'h 000200;  // +2.0000000000000000 = 2^(61+1) *  1 * atan( 1 / ( -1 + 2^61 ) )   n = 61   d_n = -1+1i 
assign v[4'b0111] [62] = 22'h 000200;  // +2.0000000000000000 = 2^(62+1) *  1 * atan( 1 / ( -1 + 2^62 ) )   n = 62   d_n = -1+1i 
assign v[4'b0111] [63] = 22'h 000200;  // +2.0000000000000000 = 2^(63+1) *  1 * atan( 1 / ( -1 + 2^63 ) )   n = 63   d_n = -1+1i 
assign v[4'b0111] [64] = 22'h 000200;  // +2.0000000000000000 = 2^(64+1) *  1 * atan( 1 / ( -1 + 2^64 ) )   n = 64   d_n = -1+1i 
assign v[4'b1000] [01] = 22'h 000000;  // +0.0000000000000000 = 2^(1+1) *  0 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = 0 
assign v[4'b1000] [02] = 22'h 000000;  // +0.0000000000000000 = 2^(2+1) *  0 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = 0 
assign v[4'b1000] [03] = 22'h 000000;  // +0.0000000000000000 = 2^(3+1) *  0 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = 0 
assign v[4'b1000] [04] = 22'h 000000;  // +0.0000000000000000 = 2^(4+1) *  0 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = 0 
assign v[4'b1000] [05] = 22'h 000000;  // +0.0000000000000000 = 2^(5+1) *  0 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = 0 
assign v[4'b1000] [06] = 22'h 000000;  // +0.0000000000000000 = 2^(6+1) *  0 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = 0 
assign v[4'b1000] [07] = 22'h 000000;  // +0.0000000000000000 = 2^(7+1) *  0 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = 0 
assign v[4'b1000] [08] = 22'h 000000;  // +0.0000000000000000 = 2^(8+1) *  0 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = 0 
assign v[4'b1000] [09] = 22'h 000000;  // +0.0000000000000000 = 2^(9+1) *  0 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = 0 
assign v[4'b1000] [10] = 22'h 000000;  // +0.0000000000000000 = 2^(10+1) *  0 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = 0 
assign v[4'b1000] [11] = 22'h 000000;  // +0.0000000000000000 = 2^(11+1) *  0 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = 0 
assign v[4'b1000] [12] = 22'h 000000;  // +0.0000000000000000 = 2^(12+1) *  0 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = 0 
assign v[4'b1000] [13] = 22'h 000000;  // +0.0000000000000000 = 2^(13+1) *  0 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = 0 
assign v[4'b1000] [14] = 22'h 000000;  // +0.0000000000000000 = 2^(14+1) *  0 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = 0 
assign v[4'b1000] [15] = 22'h 000000;  // +0.0000000000000000 = 2^(15+1) *  0 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = 0 
assign v[4'b1000] [16] = 22'h 000000;  // +0.0000000000000000 = 2^(16+1) *  0 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = 0 
assign v[4'b1000] [17] = 22'h 000000;  // +0.0000000000000000 = 2^(17+1) *  0 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = 0 
assign v[4'b1000] [18] = 22'h 000000;  // +0.0000000000000000 = 2^(18+1) *  0 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = 0 
assign v[4'b1000] [19] = 22'h 000000;  // +0.0000000000000000 = 2^(19+1) *  0 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = 0 
assign v[4'b1000] [20] = 22'h 000000;  // +0.0000000000000000 = 2^(20+1) *  0 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = 0 
assign v[4'b1000] [21] = 22'h 000000;  // +0.0000000000000000 = 2^(21+1) *  0 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = 0 
assign v[4'b1000] [22] = 22'h 000000;  // +0.0000000000000000 = 2^(22+1) *  0 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = 0 
assign v[4'b1000] [23] = 22'h 000000;  // +0.0000000000000000 = 2^(23+1) *  0 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = 0 
assign v[4'b1000] [24] = 22'h 000000;  // +0.0000000000000000 = 2^(24+1) *  0 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = 0 
assign v[4'b1000] [25] = 22'h 000000;  // +0.0000000000000000 = 2^(25+1) *  0 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = 0 
assign v[4'b1000] [26] = 22'h 000000;  // +0.0000000000000000 = 2^(26+1) *  0 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = 0 
assign v[4'b1000] [27] = 22'h 000000;  // +0.0000000000000000 = 2^(27+1) *  0 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = 0 
assign v[4'b1000] [28] = 22'h 000000;  // +0.0000000000000000 = 2^(28+1) *  0 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = 0 
assign v[4'b1000] [29] = 22'h 000000;  // +0.0000000000000000 = 2^(29+1) *  0 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = 0 
assign v[4'b1000] [30] = 22'h 000000;  // +0.0000000000000000 = 2^(30+1) *  0 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = 0 
assign v[4'b1000] [31] = 22'h 000000;  // +0.0000000000000000 = 2^(31+1) *  0 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = 0 
assign v[4'b1000] [32] = 22'h 000000;  // +0.0000000000000000 = 2^(32+1) *  0 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = 0 
assign v[4'b1000] [33] = 22'h 000000;  // +0.0000000000000000 = 2^(33+1) *  0 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = 0 
assign v[4'b1000] [34] = 22'h 000000;  // +0.0000000000000000 = 2^(34+1) *  0 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = 0 
assign v[4'b1000] [35] = 22'h 000000;  // +0.0000000000000000 = 2^(35+1) *  0 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = 0 
assign v[4'b1000] [36] = 22'h 000000;  // +0.0000000000000000 = 2^(36+1) *  0 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = 0 
assign v[4'b1000] [37] = 22'h 000000;  // +0.0000000000000000 = 2^(37+1) *  0 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = 0 
assign v[4'b1000] [38] = 22'h 000000;  // +0.0000000000000000 = 2^(38+1) *  0 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = 0 
assign v[4'b1000] [39] = 22'h 000000;  // +0.0000000000000000 = 2^(39+1) *  0 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = 0 
assign v[4'b1000] [40] = 22'h 000000;  // +0.0000000000000000 = 2^(40+1) *  0 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = 0 
assign v[4'b1000] [41] = 22'h 000000;  // +0.0000000000000000 = 2^(41+1) *  0 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = 0 
assign v[4'b1000] [42] = 22'h 000000;  // +0.0000000000000000 = 2^(42+1) *  0 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = 0 
assign v[4'b1000] [43] = 22'h 000000;  // +0.0000000000000000 = 2^(43+1) *  0 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = 0 
assign v[4'b1000] [44] = 22'h 000000;  // +0.0000000000000000 = 2^(44+1) *  0 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = 0 
assign v[4'b1000] [45] = 22'h 000000;  // +0.0000000000000000 = 2^(45+1) *  0 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = 0 
assign v[4'b1000] [46] = 22'h 000000;  // +0.0000000000000000 = 2^(46+1) *  0 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = 0 
assign v[4'b1000] [47] = 22'h 000000;  // +0.0000000000000000 = 2^(47+1) *  0 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = 0 
assign v[4'b1000] [48] = 22'h 000000;  // +0.0000000000000000 = 2^(48+1) *  0 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = 0 
assign v[4'b1000] [49] = 22'h 000000;  // +0.0000000000000000 = 2^(49+1) *  0 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = 0 
assign v[4'b1000] [50] = 22'h 000000;  // +0.0000000000000000 = 2^(50+1) *  0 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = 0 
assign v[4'b1000] [51] = 22'h 000000;  // +0.0000000000000000 = 2^(51+1) *  0 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = 0 
assign v[4'b1000] [52] = 22'h 000000;  // +0.0000000000000000 = 2^(52+1) *  0 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = 0 
assign v[4'b1000] [53] = 22'h 000000;  // +0.0000000000000000 = 2^(53+1) *  0 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = 0 
assign v[4'b1000] [54] = 22'h 000000;  // +0.0000000000000000 = 2^(54+1) *  0 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = 0 
assign v[4'b1000] [55] = 22'h 000000;  // +0.0000000000000000 = 2^(55+1) *  0 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = 0 
assign v[4'b1000] [56] = 22'h 000000;  // +0.0000000000000000 = 2^(56+1) *  0 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = 0 
assign v[4'b1000] [57] = 22'h 000000;  // +0.0000000000000000 = 2^(57+1) *  0 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = 0 
assign v[4'b1000] [58] = 22'h 000000;  // +0.0000000000000000 = 2^(58+1) *  0 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = 0 
assign v[4'b1000] [59] = 22'h 000000;  // +0.0000000000000000 = 2^(59+1) *  0 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = 0 
assign v[4'b1000] [60] = 22'h 000000;  // +0.0000000000000000 = 2^(60+1) *  0 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = 0 
assign v[4'b1000] [61] = 22'h 000000;  // +0.0000000000000000 = 2^(61+1) *  0 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = 0 
assign v[4'b1000] [62] = 22'h 000000;  // +0.0000000000000000 = 2^(62+1) *  0 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = 0 
assign v[4'b1000] [63] = 22'h 000000;  // +0.0000000000000000 = 2^(63+1) *  0 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = 0 
assign v[4'b1000] [64] = 22'h 000000;  // +0.0000000000000000 = 2^(64+1) *  0 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = 0 
assign v[4'b1001] [01] = 22'h 000000;  // +0.0000000000000000 = 2^(1+1) *  0 * atan( 1 / (  1 + 2^1 ) )   n =  1   d_n = 1 
assign v[4'b1001] [02] = 22'h 000000;  // +0.0000000000000000 = 2^(2+1) *  0 * atan( 1 / (  1 + 2^2 ) )   n =  2   d_n = 1 
assign v[4'b1001] [03] = 22'h 000000;  // +0.0000000000000000 = 2^(3+1) *  0 * atan( 1 / (  1 + 2^3 ) )   n =  3   d_n = 1 
assign v[4'b1001] [04] = 22'h 000000;  // +0.0000000000000000 = 2^(4+1) *  0 * atan( 1 / (  1 + 2^4 ) )   n =  4   d_n = 1 
assign v[4'b1001] [05] = 22'h 000000;  // +0.0000000000000000 = 2^(5+1) *  0 * atan( 1 / (  1 + 2^5 ) )   n =  5   d_n = 1 
assign v[4'b1001] [06] = 22'h 000000;  // +0.0000000000000000 = 2^(6+1) *  0 * atan( 1 / (  1 + 2^6 ) )   n =  6   d_n = 1 
assign v[4'b1001] [07] = 22'h 000000;  // +0.0000000000000000 = 2^(7+1) *  0 * atan( 1 / (  1 + 2^7 ) )   n =  7   d_n = 1 
assign v[4'b1001] [08] = 22'h 000000;  // +0.0000000000000000 = 2^(8+1) *  0 * atan( 1 / (  1 + 2^8 ) )   n =  8   d_n = 1 
assign v[4'b1001] [09] = 22'h 000000;  // +0.0000000000000000 = 2^(9+1) *  0 * atan( 1 / (  1 + 2^9 ) )   n =  9   d_n = 1 
assign v[4'b1001] [10] = 22'h 000000;  // +0.0000000000000000 = 2^(10+1) *  0 * atan( 1 / (  1 + 2^10 ) )   n = 10   d_n = 1 
assign v[4'b1001] [11] = 22'h 000000;  // +0.0000000000000000 = 2^(11+1) *  0 * atan( 1 / (  1 + 2^11 ) )   n = 11   d_n = 1 
assign v[4'b1001] [12] = 22'h 000000;  // +0.0000000000000000 = 2^(12+1) *  0 * atan( 1 / (  1 + 2^12 ) )   n = 12   d_n = 1 
assign v[4'b1001] [13] = 22'h 000000;  // +0.0000000000000000 = 2^(13+1) *  0 * atan( 1 / (  1 + 2^13 ) )   n = 13   d_n = 1 
assign v[4'b1001] [14] = 22'h 000000;  // +0.0000000000000000 = 2^(14+1) *  0 * atan( 1 / (  1 + 2^14 ) )   n = 14   d_n = 1 
assign v[4'b1001] [15] = 22'h 000000;  // +0.0000000000000000 = 2^(15+1) *  0 * atan( 1 / (  1 + 2^15 ) )   n = 15   d_n = 1 
assign v[4'b1001] [16] = 22'h 000000;  // +0.0000000000000000 = 2^(16+1) *  0 * atan( 1 / (  1 + 2^16 ) )   n = 16   d_n = 1 
assign v[4'b1001] [17] = 22'h 000000;  // +0.0000000000000000 = 2^(17+1) *  0 * atan( 1 / (  1 + 2^17 ) )   n = 17   d_n = 1 
assign v[4'b1001] [18] = 22'h 000000;  // +0.0000000000000000 = 2^(18+1) *  0 * atan( 1 / (  1 + 2^18 ) )   n = 18   d_n = 1 
assign v[4'b1001] [19] = 22'h 000000;  // +0.0000000000000000 = 2^(19+1) *  0 * atan( 1 / (  1 + 2^19 ) )   n = 19   d_n = 1 
assign v[4'b1001] [20] = 22'h 000000;  // +0.0000000000000000 = 2^(20+1) *  0 * atan( 1 / (  1 + 2^20 ) )   n = 20   d_n = 1 
assign v[4'b1001] [21] = 22'h 000000;  // +0.0000000000000000 = 2^(21+1) *  0 * atan( 1 / (  1 + 2^21 ) )   n = 21   d_n = 1 
assign v[4'b1001] [22] = 22'h 000000;  // +0.0000000000000000 = 2^(22+1) *  0 * atan( 1 / (  1 + 2^22 ) )   n = 22   d_n = 1 
assign v[4'b1001] [23] = 22'h 000000;  // +0.0000000000000000 = 2^(23+1) *  0 * atan( 1 / (  1 + 2^23 ) )   n = 23   d_n = 1 
assign v[4'b1001] [24] = 22'h 000000;  // +0.0000000000000000 = 2^(24+1) *  0 * atan( 1 / (  1 + 2^24 ) )   n = 24   d_n = 1 
assign v[4'b1001] [25] = 22'h 000000;  // +0.0000000000000000 = 2^(25+1) *  0 * atan( 1 / (  1 + 2^25 ) )   n = 25   d_n = 1 
assign v[4'b1001] [26] = 22'h 000000;  // +0.0000000000000000 = 2^(26+1) *  0 * atan( 1 / (  1 + 2^26 ) )   n = 26   d_n = 1 
assign v[4'b1001] [27] = 22'h 000000;  // +0.0000000000000000 = 2^(27+1) *  0 * atan( 1 / (  1 + 2^27 ) )   n = 27   d_n = 1 
assign v[4'b1001] [28] = 22'h 000000;  // +0.0000000000000000 = 2^(28+1) *  0 * atan( 1 / (  1 + 2^28 ) )   n = 28   d_n = 1 
assign v[4'b1001] [29] = 22'h 000000;  // +0.0000000000000000 = 2^(29+1) *  0 * atan( 1 / (  1 + 2^29 ) )   n = 29   d_n = 1 
assign v[4'b1001] [30] = 22'h 000000;  // +0.0000000000000000 = 2^(30+1) *  0 * atan( 1 / (  1 + 2^30 ) )   n = 30   d_n = 1 
assign v[4'b1001] [31] = 22'h 000000;  // +0.0000000000000000 = 2^(31+1) *  0 * atan( 1 / (  1 + 2^31 ) )   n = 31   d_n = 1 
assign v[4'b1001] [32] = 22'h 000000;  // +0.0000000000000000 = 2^(32+1) *  0 * atan( 1 / (  1 + 2^32 ) )   n = 32   d_n = 1 
assign v[4'b1001] [33] = 22'h 000000;  // +0.0000000000000000 = 2^(33+1) *  0 * atan( 1 / (  1 + 2^33 ) )   n = 33   d_n = 1 
assign v[4'b1001] [34] = 22'h 000000;  // +0.0000000000000000 = 2^(34+1) *  0 * atan( 1 / (  1 + 2^34 ) )   n = 34   d_n = 1 
assign v[4'b1001] [35] = 22'h 000000;  // +0.0000000000000000 = 2^(35+1) *  0 * atan( 1 / (  1 + 2^35 ) )   n = 35   d_n = 1 
assign v[4'b1001] [36] = 22'h 000000;  // +0.0000000000000000 = 2^(36+1) *  0 * atan( 1 / (  1 + 2^36 ) )   n = 36   d_n = 1 
assign v[4'b1001] [37] = 22'h 000000;  // +0.0000000000000000 = 2^(37+1) *  0 * atan( 1 / (  1 + 2^37 ) )   n = 37   d_n = 1 
assign v[4'b1001] [38] = 22'h 000000;  // +0.0000000000000000 = 2^(38+1) *  0 * atan( 1 / (  1 + 2^38 ) )   n = 38   d_n = 1 
assign v[4'b1001] [39] = 22'h 000000;  // +0.0000000000000000 = 2^(39+1) *  0 * atan( 1 / (  1 + 2^39 ) )   n = 39   d_n = 1 
assign v[4'b1001] [40] = 22'h 000000;  // +0.0000000000000000 = 2^(40+1) *  0 * atan( 1 / (  1 + 2^40 ) )   n = 40   d_n = 1 
assign v[4'b1001] [41] = 22'h 000000;  // +0.0000000000000000 = 2^(41+1) *  0 * atan( 1 / (  1 + 2^41 ) )   n = 41   d_n = 1 
assign v[4'b1001] [42] = 22'h 000000;  // +0.0000000000000000 = 2^(42+1) *  0 * atan( 1 / (  1 + 2^42 ) )   n = 42   d_n = 1 
assign v[4'b1001] [43] = 22'h 000000;  // +0.0000000000000000 = 2^(43+1) *  0 * atan( 1 / (  1 + 2^43 ) )   n = 43   d_n = 1 
assign v[4'b1001] [44] = 22'h 000000;  // +0.0000000000000000 = 2^(44+1) *  0 * atan( 1 / (  1 + 2^44 ) )   n = 44   d_n = 1 
assign v[4'b1001] [45] = 22'h 000000;  // +0.0000000000000000 = 2^(45+1) *  0 * atan( 1 / (  1 + 2^45 ) )   n = 45   d_n = 1 
assign v[4'b1001] [46] = 22'h 000000;  // +0.0000000000000000 = 2^(46+1) *  0 * atan( 1 / (  1 + 2^46 ) )   n = 46   d_n = 1 
assign v[4'b1001] [47] = 22'h 000000;  // +0.0000000000000000 = 2^(47+1) *  0 * atan( 1 / (  1 + 2^47 ) )   n = 47   d_n = 1 
assign v[4'b1001] [48] = 22'h 000000;  // +0.0000000000000000 = 2^(48+1) *  0 * atan( 1 / (  1 + 2^48 ) )   n = 48   d_n = 1 
assign v[4'b1001] [49] = 22'h 000000;  // +0.0000000000000000 = 2^(49+1) *  0 * atan( 1 / (  1 + 2^49 ) )   n = 49   d_n = 1 
assign v[4'b1001] [50] = 22'h 000000;  // +0.0000000000000000 = 2^(50+1) *  0 * atan( 1 / (  1 + 2^50 ) )   n = 50   d_n = 1 
assign v[4'b1001] [51] = 22'h 000000;  // +0.0000000000000000 = 2^(51+1) *  0 * atan( 1 / (  1 + 2^51 ) )   n = 51   d_n = 1 
assign v[4'b1001] [52] = 22'h 000000;  // +0.0000000000000000 = 2^(52+1) *  0 * atan( 1 / (  1 + 2^52 ) )   n = 52   d_n = 1 
assign v[4'b1001] [53] = 22'h 000000;  // +0.0000000000000000 = 2^(53+1) *  0 * atan( 1 / (  1 + 2^53 ) )   n = 53   d_n = 1 
assign v[4'b1001] [54] = 22'h 000000;  // +0.0000000000000000 = 2^(54+1) *  0 * atan( 1 / (  1 + 2^54 ) )   n = 54   d_n = 1 
assign v[4'b1001] [55] = 22'h 000000;  // +0.0000000000000000 = 2^(55+1) *  0 * atan( 1 / (  1 + 2^55 ) )   n = 55   d_n = 1 
assign v[4'b1001] [56] = 22'h 000000;  // +0.0000000000000000 = 2^(56+1) *  0 * atan( 1 / (  1 + 2^56 ) )   n = 56   d_n = 1 
assign v[4'b1001] [57] = 22'h 000000;  // +0.0000000000000000 = 2^(57+1) *  0 * atan( 1 / (  1 + 2^57 ) )   n = 57   d_n = 1 
assign v[4'b1001] [58] = 22'h 000000;  // +0.0000000000000000 = 2^(58+1) *  0 * atan( 1 / (  1 + 2^58 ) )   n = 58   d_n = 1 
assign v[4'b1001] [59] = 22'h 000000;  // +0.0000000000000000 = 2^(59+1) *  0 * atan( 1 / (  1 + 2^59 ) )   n = 59   d_n = 1 
assign v[4'b1001] [60] = 22'h 000000;  // +0.0000000000000000 = 2^(60+1) *  0 * atan( 1 / (  1 + 2^60 ) )   n = 60   d_n = 1 
assign v[4'b1001] [61] = 22'h 000000;  // +0.0000000000000000 = 2^(61+1) *  0 * atan( 1 / (  1 + 2^61 ) )   n = 61   d_n = 1 
assign v[4'b1001] [62] = 22'h 000000;  // +0.0000000000000000 = 2^(62+1) *  0 * atan( 1 / (  1 + 2^62 ) )   n = 62   d_n = 1 
assign v[4'b1001] [63] = 22'h 000000;  // +0.0000000000000000 = 2^(63+1) *  0 * atan( 1 / (  1 + 2^63 ) )   n = 63   d_n = 1 
assign v[4'b1001] [64] = 22'h 000000;  // +0.0000000000000000 = 2^(64+1) *  0 * atan( 1 / (  1 + 2^64 ) )   n = 64   d_n = 1 
assign v[4'b1010] [01] = 22'h 000000;  // +0.0000000000000000 = 2^(1+1) *  0 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = -0 
assign v[4'b1010] [02] = 22'h 000000;  // +0.0000000000000000 = 2^(2+1) *  0 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = -0 
assign v[4'b1010] [03] = 22'h 000000;  // +0.0000000000000000 = 2^(3+1) *  0 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = -0 
assign v[4'b1010] [04] = 22'h 000000;  // +0.0000000000000000 = 2^(4+1) *  0 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = -0 
assign v[4'b1010] [05] = 22'h 000000;  // +0.0000000000000000 = 2^(5+1) *  0 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = -0 
assign v[4'b1010] [06] = 22'h 000000;  // +0.0000000000000000 = 2^(6+1) *  0 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = -0 
assign v[4'b1010] [07] = 22'h 000000;  // +0.0000000000000000 = 2^(7+1) *  0 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = -0 
assign v[4'b1010] [08] = 22'h 000000;  // +0.0000000000000000 = 2^(8+1) *  0 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = -0 
assign v[4'b1010] [09] = 22'h 000000;  // +0.0000000000000000 = 2^(9+1) *  0 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = -0 
assign v[4'b1010] [10] = 22'h 000000;  // +0.0000000000000000 = 2^(10+1) *  0 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = -0 
assign v[4'b1010] [11] = 22'h 000000;  // +0.0000000000000000 = 2^(11+1) *  0 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = -0 
assign v[4'b1010] [12] = 22'h 000000;  // +0.0000000000000000 = 2^(12+1) *  0 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = -0 
assign v[4'b1010] [13] = 22'h 000000;  // +0.0000000000000000 = 2^(13+1) *  0 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = -0 
assign v[4'b1010] [14] = 22'h 000000;  // +0.0000000000000000 = 2^(14+1) *  0 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = -0 
assign v[4'b1010] [15] = 22'h 000000;  // +0.0000000000000000 = 2^(15+1) *  0 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = -0 
assign v[4'b1010] [16] = 22'h 000000;  // +0.0000000000000000 = 2^(16+1) *  0 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = -0 
assign v[4'b1010] [17] = 22'h 000000;  // +0.0000000000000000 = 2^(17+1) *  0 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = -0 
assign v[4'b1010] [18] = 22'h 000000;  // +0.0000000000000000 = 2^(18+1) *  0 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = -0 
assign v[4'b1010] [19] = 22'h 000000;  // +0.0000000000000000 = 2^(19+1) *  0 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = -0 
assign v[4'b1010] [20] = 22'h 000000;  // +0.0000000000000000 = 2^(20+1) *  0 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = -0 
assign v[4'b1010] [21] = 22'h 000000;  // +0.0000000000000000 = 2^(21+1) *  0 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = -0 
assign v[4'b1010] [22] = 22'h 000000;  // +0.0000000000000000 = 2^(22+1) *  0 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = -0 
assign v[4'b1010] [23] = 22'h 000000;  // +0.0000000000000000 = 2^(23+1) *  0 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = -0 
assign v[4'b1010] [24] = 22'h 000000;  // +0.0000000000000000 = 2^(24+1) *  0 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = -0 
assign v[4'b1010] [25] = 22'h 000000;  // +0.0000000000000000 = 2^(25+1) *  0 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = -0 
assign v[4'b1010] [26] = 22'h 000000;  // +0.0000000000000000 = 2^(26+1) *  0 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = -0 
assign v[4'b1010] [27] = 22'h 000000;  // +0.0000000000000000 = 2^(27+1) *  0 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = -0 
assign v[4'b1010] [28] = 22'h 000000;  // +0.0000000000000000 = 2^(28+1) *  0 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = -0 
assign v[4'b1010] [29] = 22'h 000000;  // +0.0000000000000000 = 2^(29+1) *  0 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = -0 
assign v[4'b1010] [30] = 22'h 000000;  // +0.0000000000000000 = 2^(30+1) *  0 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = -0 
assign v[4'b1010] [31] = 22'h 000000;  // +0.0000000000000000 = 2^(31+1) *  0 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = -0 
assign v[4'b1010] [32] = 22'h 000000;  // +0.0000000000000000 = 2^(32+1) *  0 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = -0 
assign v[4'b1010] [33] = 22'h 000000;  // +0.0000000000000000 = 2^(33+1) *  0 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = -0 
assign v[4'b1010] [34] = 22'h 000000;  // +0.0000000000000000 = 2^(34+1) *  0 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = -0 
assign v[4'b1010] [35] = 22'h 000000;  // +0.0000000000000000 = 2^(35+1) *  0 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = -0 
assign v[4'b1010] [36] = 22'h 000000;  // +0.0000000000000000 = 2^(36+1) *  0 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = -0 
assign v[4'b1010] [37] = 22'h 000000;  // +0.0000000000000000 = 2^(37+1) *  0 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = -0 
assign v[4'b1010] [38] = 22'h 000000;  // +0.0000000000000000 = 2^(38+1) *  0 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = -0 
assign v[4'b1010] [39] = 22'h 000000;  // +0.0000000000000000 = 2^(39+1) *  0 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = -0 
assign v[4'b1010] [40] = 22'h 000000;  // +0.0000000000000000 = 2^(40+1) *  0 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = -0 
assign v[4'b1010] [41] = 22'h 000000;  // +0.0000000000000000 = 2^(41+1) *  0 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = -0 
assign v[4'b1010] [42] = 22'h 000000;  // +0.0000000000000000 = 2^(42+1) *  0 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = -0 
assign v[4'b1010] [43] = 22'h 000000;  // +0.0000000000000000 = 2^(43+1) *  0 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = -0 
assign v[4'b1010] [44] = 22'h 000000;  // +0.0000000000000000 = 2^(44+1) *  0 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = -0 
assign v[4'b1010] [45] = 22'h 000000;  // +0.0000000000000000 = 2^(45+1) *  0 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = -0 
assign v[4'b1010] [46] = 22'h 000000;  // +0.0000000000000000 = 2^(46+1) *  0 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = -0 
assign v[4'b1010] [47] = 22'h 000000;  // +0.0000000000000000 = 2^(47+1) *  0 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = -0 
assign v[4'b1010] [48] = 22'h 000000;  // +0.0000000000000000 = 2^(48+1) *  0 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = -0 
assign v[4'b1010] [49] = 22'h 000000;  // +0.0000000000000000 = 2^(49+1) *  0 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = -0 
assign v[4'b1010] [50] = 22'h 000000;  // +0.0000000000000000 = 2^(50+1) *  0 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = -0 
assign v[4'b1010] [51] = 22'h 000000;  // +0.0000000000000000 = 2^(51+1) *  0 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = -0 
assign v[4'b1010] [52] = 22'h 000000;  // +0.0000000000000000 = 2^(52+1) *  0 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = -0 
assign v[4'b1010] [53] = 22'h 000000;  // +0.0000000000000000 = 2^(53+1) *  0 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = -0 
assign v[4'b1010] [54] = 22'h 000000;  // +0.0000000000000000 = 2^(54+1) *  0 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = -0 
assign v[4'b1010] [55] = 22'h 000000;  // +0.0000000000000000 = 2^(55+1) *  0 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = -0 
assign v[4'b1010] [56] = 22'h 000000;  // +0.0000000000000000 = 2^(56+1) *  0 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = -0 
assign v[4'b1010] [57] = 22'h 000000;  // +0.0000000000000000 = 2^(57+1) *  0 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = -0 
assign v[4'b1010] [58] = 22'h 000000;  // +0.0000000000000000 = 2^(58+1) *  0 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = -0 
assign v[4'b1010] [59] = 22'h 000000;  // +0.0000000000000000 = 2^(59+1) *  0 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = -0 
assign v[4'b1010] [60] = 22'h 000000;  // +0.0000000000000000 = 2^(60+1) *  0 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = -0 
assign v[4'b1010] [61] = 22'h 000000;  // +0.0000000000000000 = 2^(61+1) *  0 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = -0 
assign v[4'b1010] [62] = 22'h 000000;  // +0.0000000000000000 = 2^(62+1) *  0 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = -0 
assign v[4'b1010] [63] = 22'h 000000;  // +0.0000000000000000 = 2^(63+1) *  0 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = -0 
assign v[4'b1010] [64] = 22'h 000000;  // +0.0000000000000000 = 2^(64+1) *  0 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = -0 
assign v[4'b1011] [01] = 22'h 000000;  // -0.0000000000000000 = 2^(1+1) *  0 * atan( 1 / ( -1 + 2^1 ) )   n =  1   d_n = -1 
assign v[4'b1011] [02] = 22'h 000000;  // -0.0000000000000000 = 2^(2+1) *  0 * atan( 1 / ( -1 + 2^2 ) )   n =  2   d_n = -1 
assign v[4'b1011] [03] = 22'h 000000;  // -0.0000000000000000 = 2^(3+1) *  0 * atan( 1 / ( -1 + 2^3 ) )   n =  3   d_n = -1 
assign v[4'b1011] [04] = 22'h 000000;  // -0.0000000000000000 = 2^(4+1) *  0 * atan( 1 / ( -1 + 2^4 ) )   n =  4   d_n = -1 
assign v[4'b1011] [05] = 22'h 000000;  // -0.0000000000000000 = 2^(5+1) *  0 * atan( 1 / ( -1 + 2^5 ) )   n =  5   d_n = -1 
assign v[4'b1011] [06] = 22'h 000000;  // -0.0000000000000000 = 2^(6+1) *  0 * atan( 1 / ( -1 + 2^6 ) )   n =  6   d_n = -1 
assign v[4'b1011] [07] = 22'h 000000;  // -0.0000000000000000 = 2^(7+1) *  0 * atan( 1 / ( -1 + 2^7 ) )   n =  7   d_n = -1 
assign v[4'b1011] [08] = 22'h 000000;  // -0.0000000000000000 = 2^(8+1) *  0 * atan( 1 / ( -1 + 2^8 ) )   n =  8   d_n = -1 
assign v[4'b1011] [09] = 22'h 000000;  // -0.0000000000000000 = 2^(9+1) *  0 * atan( 1 / ( -1 + 2^9 ) )   n =  9   d_n = -1 
assign v[4'b1011] [10] = 22'h 000000;  // -0.0000000000000000 = 2^(10+1) *  0 * atan( 1 / ( -1 + 2^10 ) )   n = 10   d_n = -1 
assign v[4'b1011] [11] = 22'h 000000;  // -0.0000000000000000 = 2^(11+1) *  0 * atan( 1 / ( -1 + 2^11 ) )   n = 11   d_n = -1 
assign v[4'b1011] [12] = 22'h 000000;  // -0.0000000000000000 = 2^(12+1) *  0 * atan( 1 / ( -1 + 2^12 ) )   n = 12   d_n = -1 
assign v[4'b1011] [13] = 22'h 000000;  // -0.0000000000000000 = 2^(13+1) *  0 * atan( 1 / ( -1 + 2^13 ) )   n = 13   d_n = -1 
assign v[4'b1011] [14] = 22'h 000000;  // -0.0000000000000000 = 2^(14+1) *  0 * atan( 1 / ( -1 + 2^14 ) )   n = 14   d_n = -1 
assign v[4'b1011] [15] = 22'h 000000;  // -0.0000000000000000 = 2^(15+1) *  0 * atan( 1 / ( -1 + 2^15 ) )   n = 15   d_n = -1 
assign v[4'b1011] [16] = 22'h 000000;  // -0.0000000000000000 = 2^(16+1) *  0 * atan( 1 / ( -1 + 2^16 ) )   n = 16   d_n = -1 
assign v[4'b1011] [17] = 22'h 000000;  // -0.0000000000000000 = 2^(17+1) *  0 * atan( 1 / ( -1 + 2^17 ) )   n = 17   d_n = -1 
assign v[4'b1011] [18] = 22'h 000000;  // -0.0000000000000000 = 2^(18+1) *  0 * atan( 1 / ( -1 + 2^18 ) )   n = 18   d_n = -1 
assign v[4'b1011] [19] = 22'h 000000;  // -0.0000000000000000 = 2^(19+1) *  0 * atan( 1 / ( -1 + 2^19 ) )   n = 19   d_n = -1 
assign v[4'b1011] [20] = 22'h 000000;  // -0.0000000000000000 = 2^(20+1) *  0 * atan( 1 / ( -1 + 2^20 ) )   n = 20   d_n = -1 
assign v[4'b1011] [21] = 22'h 000000;  // -0.0000000000000000 = 2^(21+1) *  0 * atan( 1 / ( -1 + 2^21 ) )   n = 21   d_n = -1 
assign v[4'b1011] [22] = 22'h 000000;  // -0.0000000000000000 = 2^(22+1) *  0 * atan( 1 / ( -1 + 2^22 ) )   n = 22   d_n = -1 
assign v[4'b1011] [23] = 22'h 000000;  // -0.0000000000000000 = 2^(23+1) *  0 * atan( 1 / ( -1 + 2^23 ) )   n = 23   d_n = -1 
assign v[4'b1011] [24] = 22'h 000000;  // -0.0000000000000000 = 2^(24+1) *  0 * atan( 1 / ( -1 + 2^24 ) )   n = 24   d_n = -1 
assign v[4'b1011] [25] = 22'h 000000;  // -0.0000000000000000 = 2^(25+1) *  0 * atan( 1 / ( -1 + 2^25 ) )   n = 25   d_n = -1 
assign v[4'b1011] [26] = 22'h 000000;  // -0.0000000000000000 = 2^(26+1) *  0 * atan( 1 / ( -1 + 2^26 ) )   n = 26   d_n = -1 
assign v[4'b1011] [27] = 22'h 000000;  // -0.0000000000000000 = 2^(27+1) *  0 * atan( 1 / ( -1 + 2^27 ) )   n = 27   d_n = -1 
assign v[4'b1011] [28] = 22'h 000000;  // -0.0000000000000000 = 2^(28+1) *  0 * atan( 1 / ( -1 + 2^28 ) )   n = 28   d_n = -1 
assign v[4'b1011] [29] = 22'h 000000;  // -0.0000000000000000 = 2^(29+1) *  0 * atan( 1 / ( -1 + 2^29 ) )   n = 29   d_n = -1 
assign v[4'b1011] [30] = 22'h 000000;  // -0.0000000000000000 = 2^(30+1) *  0 * atan( 1 / ( -1 + 2^30 ) )   n = 30   d_n = -1 
assign v[4'b1011] [31] = 22'h 000000;  // -0.0000000000000000 = 2^(31+1) *  0 * atan( 1 / ( -1 + 2^31 ) )   n = 31   d_n = -1 
assign v[4'b1011] [32] = 22'h 000000;  // -0.0000000000000000 = 2^(32+1) *  0 * atan( 1 / ( -1 + 2^32 ) )   n = 32   d_n = -1 
assign v[4'b1011] [33] = 22'h 000000;  // -0.0000000000000000 = 2^(33+1) *  0 * atan( 1 / ( -1 + 2^33 ) )   n = 33   d_n = -1 
assign v[4'b1011] [34] = 22'h 000000;  // -0.0000000000000000 = 2^(34+1) *  0 * atan( 1 / ( -1 + 2^34 ) )   n = 34   d_n = -1 
assign v[4'b1011] [35] = 22'h 000000;  // -0.0000000000000000 = 2^(35+1) *  0 * atan( 1 / ( -1 + 2^35 ) )   n = 35   d_n = -1 
assign v[4'b1011] [36] = 22'h 000000;  // -0.0000000000000000 = 2^(36+1) *  0 * atan( 1 / ( -1 + 2^36 ) )   n = 36   d_n = -1 
assign v[4'b1011] [37] = 22'h 000000;  // -0.0000000000000000 = 2^(37+1) *  0 * atan( 1 / ( -1 + 2^37 ) )   n = 37   d_n = -1 
assign v[4'b1011] [38] = 22'h 000000;  // -0.0000000000000000 = 2^(38+1) *  0 * atan( 1 / ( -1 + 2^38 ) )   n = 38   d_n = -1 
assign v[4'b1011] [39] = 22'h 000000;  // -0.0000000000000000 = 2^(39+1) *  0 * atan( 1 / ( -1 + 2^39 ) )   n = 39   d_n = -1 
assign v[4'b1011] [40] = 22'h 000000;  // -0.0000000000000000 = 2^(40+1) *  0 * atan( 1 / ( -1 + 2^40 ) )   n = 40   d_n = -1 
assign v[4'b1011] [41] = 22'h 000000;  // -0.0000000000000000 = 2^(41+1) *  0 * atan( 1 / ( -1 + 2^41 ) )   n = 41   d_n = -1 
assign v[4'b1011] [42] = 22'h 000000;  // -0.0000000000000000 = 2^(42+1) *  0 * atan( 1 / ( -1 + 2^42 ) )   n = 42   d_n = -1 
assign v[4'b1011] [43] = 22'h 000000;  // -0.0000000000000000 = 2^(43+1) *  0 * atan( 1 / ( -1 + 2^43 ) )   n = 43   d_n = -1 
assign v[4'b1011] [44] = 22'h 000000;  // -0.0000000000000000 = 2^(44+1) *  0 * atan( 1 / ( -1 + 2^44 ) )   n = 44   d_n = -1 
assign v[4'b1011] [45] = 22'h 000000;  // -0.0000000000000000 = 2^(45+1) *  0 * atan( 1 / ( -1 + 2^45 ) )   n = 45   d_n = -1 
assign v[4'b1011] [46] = 22'h 000000;  // -0.0000000000000000 = 2^(46+1) *  0 * atan( 1 / ( -1 + 2^46 ) )   n = 46   d_n = -1 
assign v[4'b1011] [47] = 22'h 000000;  // -0.0000000000000000 = 2^(47+1) *  0 * atan( 1 / ( -1 + 2^47 ) )   n = 47   d_n = -1 
assign v[4'b1011] [48] = 22'h 000000;  // -0.0000000000000000 = 2^(48+1) *  0 * atan( 1 / ( -1 + 2^48 ) )   n = 48   d_n = -1 
assign v[4'b1011] [49] = 22'h 000000;  // -0.0000000000000000 = 2^(49+1) *  0 * atan( 1 / ( -1 + 2^49 ) )   n = 49   d_n = -1 
assign v[4'b1011] [50] = 22'h 000000;  // -0.0000000000000000 = 2^(50+1) *  0 * atan( 1 / ( -1 + 2^50 ) )   n = 50   d_n = -1 
assign v[4'b1011] [51] = 22'h 000000;  // -0.0000000000000000 = 2^(51+1) *  0 * atan( 1 / ( -1 + 2^51 ) )   n = 51   d_n = -1 
assign v[4'b1011] [52] = 22'h 000000;  // -0.0000000000000000 = 2^(52+1) *  0 * atan( 1 / ( -1 + 2^52 ) )   n = 52   d_n = -1 
assign v[4'b1011] [53] = 22'h 000000;  // -0.0000000000000000 = 2^(53+1) *  0 * atan( 1 / ( -1 + 2^53 ) )   n = 53   d_n = -1 
assign v[4'b1011] [54] = 22'h 000000;  // -0.0000000000000000 = 2^(54+1) *  0 * atan( 1 / ( -1 + 2^54 ) )   n = 54   d_n = -1 
assign v[4'b1011] [55] = 22'h 000000;  // -0.0000000000000000 = 2^(55+1) *  0 * atan( 1 / ( -1 + 2^55 ) )   n = 55   d_n = -1 
assign v[4'b1011] [56] = 22'h 000000;  // -0.0000000000000000 = 2^(56+1) *  0 * atan( 1 / ( -1 + 2^56 ) )   n = 56   d_n = -1 
assign v[4'b1011] [57] = 22'h 000000;  // -0.0000000000000000 = 2^(57+1) *  0 * atan( 1 / ( -1 + 2^57 ) )   n = 57   d_n = -1 
assign v[4'b1011] [58] = 22'h 000000;  // -0.0000000000000000 = 2^(58+1) *  0 * atan( 1 / ( -1 + 2^58 ) )   n = 58   d_n = -1 
assign v[4'b1011] [59] = 22'h 000000;  // -0.0000000000000000 = 2^(59+1) *  0 * atan( 1 / ( -1 + 2^59 ) )   n = 59   d_n = -1 
assign v[4'b1011] [60] = 22'h 000000;  // -0.0000000000000000 = 2^(60+1) *  0 * atan( 1 / ( -1 + 2^60 ) )   n = 60   d_n = -1 
assign v[4'b1011] [61] = 22'h 000000;  // -0.0000000000000000 = 2^(61+1) *  0 * atan( 1 / ( -1 + 2^61 ) )   n = 61   d_n = -1 
assign v[4'b1011] [62] = 22'h 000000;  // -0.0000000000000000 = 2^(62+1) *  0 * atan( 1 / ( -1 + 2^62 ) )   n = 62   d_n = -1 
assign v[4'b1011] [63] = 22'h 000000;  // -0.0000000000000000 = 2^(63+1) *  0 * atan( 1 / ( -1 + 2^63 ) )   n = 63   d_n = -1 
assign v[4'b1011] [64] = 22'h 000000;  // -0.0000000000000000 = 2^(64+1) *  0 * atan( 1 / ( -1 + 2^64 ) )   n = 64   d_n = -1 
assign v[4'b1100] [01] = 22'h 3FFE25;  // -1.8545904360032244 = 2^(1+1) * -1 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = -0-1i 
assign v[4'b1100] [02] = 22'h 3FFE0A;  // -1.9598293050149131 = 2^(2+1) * -1 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = -0-1i 
assign v[4'b1100] [03] = 22'h 3FFE02;  // -1.9896799127481830 = 2^(3+1) * -1 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = -0-1i 
assign v[4'b1100] [04] = 22'h 3FFE00;  // -1.9974019198706352 = 2^(4+1) * -1 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = -0-1i 
assign v[4'b1100] [05] = 22'h 3FFE00;  // -1.9993493395371698 = 2^(5+1) * -1 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = -0-1i 
assign v[4'b1100] [06] = 22'h 3FFE00;  // -1.9998372634210344 = 2^(6+1) * -1 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = -0-1i 
assign v[4'b1100] [07] = 22'h 3FFE00;  // -1.9999593113858845 = 2^(7+1) * -1 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = -0-1i 
assign v[4'b1100] [08] = 22'h 3FFE00;  // -1.9999898275670895 = 2^(8+1) * -1 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = -0-1i 
assign v[4'b1100] [09] = 22'h 3FFE00;  // -1.9999974568743104 = 2^(9+1) * -1 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = -0-1i 
assign v[4'b1100] [10] = 22'h 3FFE00;  // -1.9999993642174863 = 2^(10+1) * -1 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = -0-1i 
assign v[4'b1100] [11] = 22'h 3FFE00;  // -1.9999998410543034 = 2^(11+1) * -1 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = -0-1i 
assign v[4'b1100] [12] = 22'h 3FFE00;  // -1.9999999602635716 = 2^(12+1) * -1 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = -0-1i 
assign v[4'b1100] [13] = 22'h 3FFE00;  // -1.9999999900658927 = 2^(13+1) * -1 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = -0-1i 
assign v[4'b1100] [14] = 22'h 3FFE00;  // -1.9999999975164731 = 2^(14+1) * -1 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = -0-1i 
assign v[4'b1100] [15] = 22'h 3FFE00;  // -1.9999999993791182 = 2^(15+1) * -1 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = -0-1i 
assign v[4'b1100] [16] = 22'h 3FFE00;  // -1.9999999998447795 = 2^(16+1) * -1 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = -0-1i 
assign v[4'b1100] [17] = 22'h 3FFE00;  // -1.9999999999611948 = 2^(17+1) * -1 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = -0-1i 
assign v[4'b1100] [18] = 22'h 3FFE00;  // -1.9999999999902986 = 2^(18+1) * -1 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = -0-1i 
assign v[4'b1100] [19] = 22'h 3FFE00;  // -1.9999999999975746 = 2^(19+1) * -1 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = -0-1i 
assign v[4'b1100] [20] = 22'h 3FFE00;  // -1.9999999999993936 = 2^(20+1) * -1 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = -0-1i 
assign v[4'b1100] [21] = 22'h 3FFE00;  // -1.9999999999998483 = 2^(21+1) * -1 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = -0-1i 
assign v[4'b1100] [22] = 22'h 3FFE00;  // -1.9999999999999620 = 2^(22+1) * -1 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = -0-1i 
assign v[4'b1100] [23] = 22'h 3FFE00;  // -1.9999999999999905 = 2^(23+1) * -1 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = -0-1i 
assign v[4'b1100] [24] = 22'h 3FFE00;  // -1.9999999999999976 = 2^(24+1) * -1 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = -0-1i 
assign v[4'b1100] [25] = 22'h 3FFE00;  // -1.9999999999999993 = 2^(25+1) * -1 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = -0-1i 
assign v[4'b1100] [26] = 22'h 3FFE00;  // -1.9999999999999998 = 2^(26+1) * -1 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = -0-1i 
assign v[4'b1100] [27] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(27+1) * -1 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = -0-1i 
assign v[4'b1100] [28] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(28+1) * -1 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = -0-1i 
assign v[4'b1100] [29] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(29+1) * -1 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = -0-1i 
assign v[4'b1100] [30] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(30+1) * -1 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = -0-1i 
assign v[4'b1100] [31] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(31+1) * -1 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = -0-1i 
assign v[4'b1100] [32] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(32+1) * -1 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = -0-1i 
assign v[4'b1100] [33] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(33+1) * -1 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = -0-1i 
assign v[4'b1100] [34] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(34+1) * -1 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = -0-1i 
assign v[4'b1100] [35] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(35+1) * -1 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = -0-1i 
assign v[4'b1100] [36] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(36+1) * -1 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = -0-1i 
assign v[4'b1100] [37] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(37+1) * -1 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = -0-1i 
assign v[4'b1100] [38] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(38+1) * -1 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = -0-1i 
assign v[4'b1100] [39] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(39+1) * -1 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = -0-1i 
assign v[4'b1100] [40] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(40+1) * -1 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = -0-1i 
assign v[4'b1100] [41] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(41+1) * -1 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = -0-1i 
assign v[4'b1100] [42] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(42+1) * -1 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = -0-1i 
assign v[4'b1100] [43] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(43+1) * -1 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = -0-1i 
assign v[4'b1100] [44] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(44+1) * -1 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = -0-1i 
assign v[4'b1100] [45] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(45+1) * -1 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = -0-1i 
assign v[4'b1100] [46] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(46+1) * -1 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = -0-1i 
assign v[4'b1100] [47] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(47+1) * -1 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = -0-1i 
assign v[4'b1100] [48] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(48+1) * -1 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = -0-1i 
assign v[4'b1100] [49] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(49+1) * -1 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = -0-1i 
assign v[4'b1100] [50] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(50+1) * -1 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = -0-1i 
assign v[4'b1100] [51] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(51+1) * -1 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = -0-1i 
assign v[4'b1100] [52] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(52+1) * -1 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = -0-1i 
assign v[4'b1100] [53] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(53+1) * -1 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = -0-1i 
assign v[4'b1100] [54] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(54+1) * -1 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = -0-1i 
assign v[4'b1100] [55] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(55+1) * -1 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = -0-1i 
assign v[4'b1100] [56] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(56+1) * -1 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = -0-1i 
assign v[4'b1100] [57] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(57+1) * -1 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = -0-1i 
assign v[4'b1100] [58] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(58+1) * -1 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = -0-1i 
assign v[4'b1100] [59] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(59+1) * -1 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = -0-1i 
assign v[4'b1100] [60] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(60+1) * -1 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = -0-1i 
assign v[4'b1100] [61] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(61+1) * -1 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = -0-1i 
assign v[4'b1100] [62] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(62+1) * -1 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = -0-1i 
assign v[4'b1100] [63] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(63+1) * -1 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = -0-1i 
assign v[4'b1100] [64] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(64+1) * -1 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = -0-1i 
assign v[4'b1101] [01] = 22'h 3FFEB6;  // -1.2870022175865687 = 2^(1+1) * -1 * atan( 1 / (  1 + 2^1 ) )   n =  1   d_n = 1-1i 
assign v[4'b1101] [02] = 22'h 3FFE6B;  // -1.5791644787990460 = 2^(2+1) * -1 * atan( 1 / (  1 + 2^2 ) )   n =  2   d_n = 1-1i 
assign v[4'b1101] [03] = 22'h 3FFE3A;  // -1.7705155387823304 = 2^(3+1) * -1 * atan( 1 / (  1 + 2^3 ) )   n =  3   d_n = 1-1i 
assign v[4'b1101] [04] = 22'h 3FFE1E;  // -1.8801863269031263 = 2^(4+1) * -1 * atan( 1 / (  1 + 2^4 ) )   n =  4   d_n = 1-1i 
assign v[4'b1101] [05] = 22'h 3FFE0F;  // -1.9388006348016065 = 2^(5+1) * -1 * atan( 1 / (  1 + 2^5 ) )   n =  5   d_n = 1-1i 
assign v[4'b1101] [06] = 22'h 3FFE07;  // -1.9690754279161793 = 2^(6+1) * -1 * atan( 1 / (  1 + 2^6 ) )   n =  6   d_n = 1-1i 
assign v[4'b1101] [07] = 22'h 3FFE03;  // -1.9844563743249595 = 2^(7+1) * -1 * atan( 1 / (  1 + 2^7 ) )   n =  7   d_n = 1-1i 
assign v[4'b1101] [08] = 22'h 3FFE01;  // -1.9922078446819715 = 2^(8+1) * -1 * atan( 1 / (  1 + 2^8 ) )   n =  8   d_n = 1-1i 
assign v[4'b1101] [09] = 22'h 3FFE00;  // -1.9960988362398133 = 2^(9+1) * -1 * atan( 1 / (  1 + 2^9 ) )   n =  9   d_n = 1-1i 
assign v[4'b1101] [10] = 22'h 3FFE00;  // -1.9980481465643023 = 2^(10+1) * -1 * atan( 1 / (  1 + 2^10 ) )   n = 10   d_n = 1-1i 
assign v[4'b1101] [11] = 22'h 3FFE00;  // -1.9990237553913479 = 2^(11+1) * -1 * atan( 1 / (  1 + 2^11 ) )   n = 11   d_n = 1-1i 
assign v[4'b1101] [12] = 22'h 3FFE00;  // -1.9995117982228541 = 2^(12+1) * -1 * atan( 1 / (  1 + 2^12 ) )   n = 12   d_n = 1-1i 
assign v[4'b1101] [13] = 22'h 3FFE00;  // -1.9997558792432146 = 2^(13+1) * -1 * atan( 1 / (  1 + 2^13 ) )   n = 13   d_n = 1-1i 
assign v[4'b1101] [14] = 22'h 3FFE00;  // -1.9998779346545537 = 2^(14+1) * -1 * atan( 1 / (  1 + 2^14 ) )   n = 14   d_n = 1-1i 
assign v[4'b1101] [15] = 22'h 3FFE00;  // -1.9999389660855134 = 2^(15+1) * -1 * atan( 1 / (  1 + 2^15 ) )   n = 15   d_n = 1-1i 
assign v[4'b1101] [16] = 22'h 3FFE00;  // -1.9999694827323158 = 2^(16+1) * -1 * atan( 1 / (  1 + 2^16 ) )   n = 16   d_n = 1-1i 
assign v[4'b1101] [17] = 22'h 3FFE00;  // -1.9999847412885476 = 2^(17+1) * -1 * atan( 1 / (  1 + 2^17 ) )   n = 17   d_n = 1-1i 
assign v[4'b1101] [18] = 22'h 3FFE00;  // -1.9999923706248712 = 2^(18+1) * -1 * atan( 1 / (  1 + 2^18 ) )   n = 18   d_n = 1-1i 
assign v[4'b1101] [19] = 22'h 3FFE00;  // -1.9999961853075849 = 2^(19+1) * -1 * atan( 1 / (  1 + 2^19 ) )   n = 19   d_n = 1-1i 
assign v[4'b1101] [20] = 22'h 3FFE00;  // -1.9999980926525798 = 2^(20+1) * -1 * atan( 1 / (  1 + 2^20 ) )   n = 20   d_n = 1-1i 
assign v[4'b1101] [21] = 22'h 3FFE00;  // -1.9999990463259867 = 2^(21+1) * -1 * atan( 1 / (  1 + 2^21 ) )   n = 21   d_n = 1-1i 
assign v[4'b1101] [22] = 22'h 3FFE00;  // -1.9999995231629175 = 2^(22+1) * -1 * atan( 1 / (  1 + 2^22 ) )   n = 22   d_n = 1-1i 
assign v[4'b1101] [23] = 22'h 3FFE00;  // -1.9999997615814398 = 2^(23+1) * -1 * atan( 1 / (  1 + 2^23 ) )   n = 23   d_n = 1-1i 
assign v[4'b1101] [24] = 22'h 3FFE00;  // -1.9999998807907151 = 2^(24+1) * -1 * atan( 1 / (  1 + 2^24 ) )   n = 24   d_n = 1-1i 
assign v[4'b1101] [25] = 22'h 3FFE00;  // -1.9999999403953563 = 2^(25+1) * -1 * atan( 1 / (  1 + 2^25 ) )   n = 25   d_n = 1-1i 
assign v[4'b1101] [26] = 22'h 3FFE00;  // -1.9999999701976778 = 2^(26+1) * -1 * atan( 1 / (  1 + 2^26 ) )   n = 26   d_n = 1-1i 
assign v[4'b1101] [27] = 22'h 3FFE00;  // -1.9999999850988388 = 2^(27+1) * -1 * atan( 1 / (  1 + 2^27 ) )   n = 27   d_n = 1-1i 
assign v[4'b1101] [28] = 22'h 3FFE00;  // -1.9999999925494194 = 2^(28+1) * -1 * atan( 1 / (  1 + 2^28 ) )   n = 28   d_n = 1-1i 
assign v[4'b1101] [29] = 22'h 3FFE00;  // -1.9999999962747097 = 2^(29+1) * -1 * atan( 1 / (  1 + 2^29 ) )   n = 29   d_n = 1-1i 
assign v[4'b1101] [30] = 22'h 3FFE00;  // -1.9999999981373549 = 2^(30+1) * -1 * atan( 1 / (  1 + 2^30 ) )   n = 30   d_n = 1-1i 
assign v[4'b1101] [31] = 22'h 3FFE00;  // -1.9999999990686774 = 2^(31+1) * -1 * atan( 1 / (  1 + 2^31 ) )   n = 31   d_n = 1-1i 
assign v[4'b1101] [32] = 22'h 3FFE00;  // -1.9999999995343387 = 2^(32+1) * -1 * atan( 1 / (  1 + 2^32 ) )   n = 32   d_n = 1-1i 
assign v[4'b1101] [33] = 22'h 3FFE00;  // -1.9999999997671694 = 2^(33+1) * -1 * atan( 1 / (  1 + 2^33 ) )   n = 33   d_n = 1-1i 
assign v[4'b1101] [34] = 22'h 3FFE00;  // -1.9999999998835847 = 2^(34+1) * -1 * atan( 1 / (  1 + 2^34 ) )   n = 34   d_n = 1-1i 
assign v[4'b1101] [35] = 22'h 3FFE00;  // -1.9999999999417923 = 2^(35+1) * -1 * atan( 1 / (  1 + 2^35 ) )   n = 35   d_n = 1-1i 
assign v[4'b1101] [36] = 22'h 3FFE00;  // -1.9999999999708962 = 2^(36+1) * -1 * atan( 1 / (  1 + 2^36 ) )   n = 36   d_n = 1-1i 
assign v[4'b1101] [37] = 22'h 3FFE00;  // -1.9999999999854481 = 2^(37+1) * -1 * atan( 1 / (  1 + 2^37 ) )   n = 37   d_n = 1-1i 
assign v[4'b1101] [38] = 22'h 3FFE00;  // -1.9999999999927240 = 2^(38+1) * -1 * atan( 1 / (  1 + 2^38 ) )   n = 38   d_n = 1-1i 
assign v[4'b1101] [39] = 22'h 3FFE00;  // -1.9999999999963620 = 2^(39+1) * -1 * atan( 1 / (  1 + 2^39 ) )   n = 39   d_n = 1-1i 
assign v[4'b1101] [40] = 22'h 3FFE00;  // -1.9999999999981810 = 2^(40+1) * -1 * atan( 1 / (  1 + 2^40 ) )   n = 40   d_n = 1-1i 
assign v[4'b1101] [41] = 22'h 3FFE00;  // -1.9999999999990905 = 2^(41+1) * -1 * atan( 1 / (  1 + 2^41 ) )   n = 41   d_n = 1-1i 
assign v[4'b1101] [42] = 22'h 3FFE00;  // -1.9999999999995453 = 2^(42+1) * -1 * atan( 1 / (  1 + 2^42 ) )   n = 42   d_n = 1-1i 
assign v[4'b1101] [43] = 22'h 3FFE00;  // -1.9999999999997726 = 2^(43+1) * -1 * atan( 1 / (  1 + 2^43 ) )   n = 43   d_n = 1-1i 
assign v[4'b1101] [44] = 22'h 3FFE00;  // -1.9999999999998863 = 2^(44+1) * -1 * atan( 1 / (  1 + 2^44 ) )   n = 44   d_n = 1-1i 
assign v[4'b1101] [45] = 22'h 3FFE00;  // -1.9999999999999432 = 2^(45+1) * -1 * atan( 1 / (  1 + 2^45 ) )   n = 45   d_n = 1-1i 
assign v[4'b1101] [46] = 22'h 3FFE00;  // -1.9999999999999716 = 2^(46+1) * -1 * atan( 1 / (  1 + 2^46 ) )   n = 46   d_n = 1-1i 
assign v[4'b1101] [47] = 22'h 3FFE00;  // -1.9999999999999858 = 2^(47+1) * -1 * atan( 1 / (  1 + 2^47 ) )   n = 47   d_n = 1-1i 
assign v[4'b1101] [48] = 22'h 3FFE00;  // -1.9999999999999929 = 2^(48+1) * -1 * atan( 1 / (  1 + 2^48 ) )   n = 48   d_n = 1-1i 
assign v[4'b1101] [49] = 22'h 3FFE00;  // -1.9999999999999964 = 2^(49+1) * -1 * atan( 1 / (  1 + 2^49 ) )   n = 49   d_n = 1-1i 
assign v[4'b1101] [50] = 22'h 3FFE00;  // -1.9999999999999982 = 2^(50+1) * -1 * atan( 1 / (  1 + 2^50 ) )   n = 50   d_n = 1-1i 
assign v[4'b1101] [51] = 22'h 3FFE00;  // -1.9999999999999991 = 2^(51+1) * -1 * atan( 1 / (  1 + 2^51 ) )   n = 51   d_n = 1-1i 
assign v[4'b1101] [52] = 22'h 3FFE00;  // -1.9999999999999996 = 2^(52+1) * -1 * atan( 1 / (  1 + 2^52 ) )   n = 52   d_n = 1-1i 
assign v[4'b1101] [53] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(53+1) * -1 * atan( 1 / (  1 + 2^53 ) )   n = 53   d_n = 1-1i 
assign v[4'b1101] [54] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(54+1) * -1 * atan( 1 / (  1 + 2^54 ) )   n = 54   d_n = 1-1i 
assign v[4'b1101] [55] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(55+1) * -1 * atan( 1 / (  1 + 2^55 ) )   n = 55   d_n = 1-1i 
assign v[4'b1101] [56] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(56+1) * -1 * atan( 1 / (  1 + 2^56 ) )   n = 56   d_n = 1-1i 
assign v[4'b1101] [57] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(57+1) * -1 * atan( 1 / (  1 + 2^57 ) )   n = 57   d_n = 1-1i 
assign v[4'b1101] [58] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(58+1) * -1 * atan( 1 / (  1 + 2^58 ) )   n = 58   d_n = 1-1i 
assign v[4'b1101] [59] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(59+1) * -1 * atan( 1 / (  1 + 2^59 ) )   n = 59   d_n = 1-1i 
assign v[4'b1101] [60] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(60+1) * -1 * atan( 1 / (  1 + 2^60 ) )   n = 60   d_n = 1-1i 
assign v[4'b1101] [61] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(61+1) * -1 * atan( 1 / (  1 + 2^61 ) )   n = 61   d_n = 1-1i 
assign v[4'b1101] [62] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(62+1) * -1 * atan( 1 / (  1 + 2^62 ) )   n = 62   d_n = 1-1i 
assign v[4'b1101] [63] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(63+1) * -1 * atan( 1 / (  1 + 2^63 ) )   n = 63   d_n = 1-1i 
assign v[4'b1101] [64] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(64+1) * -1 * atan( 1 / (  1 + 2^64 ) )   n = 64   d_n = 1-1i 
assign v[4'b1110] [01] = 22'h 3FFE25;  // -1.8545904360032244 = 2^(1+1) * -1 * atan( 1 / (  0 + 2^1 ) )   n =  1   d_n = -0-1i 
assign v[4'b1110] [02] = 22'h 3FFE0A;  // -1.9598293050149131 = 2^(2+1) * -1 * atan( 1 / (  0 + 2^2 ) )   n =  2   d_n = -0-1i 
assign v[4'b1110] [03] = 22'h 3FFE02;  // -1.9896799127481830 = 2^(3+1) * -1 * atan( 1 / (  0 + 2^3 ) )   n =  3   d_n = -0-1i 
assign v[4'b1110] [04] = 22'h 3FFE00;  // -1.9974019198706352 = 2^(4+1) * -1 * atan( 1 / (  0 + 2^4 ) )   n =  4   d_n = -0-1i 
assign v[4'b1110] [05] = 22'h 3FFE00;  // -1.9993493395371698 = 2^(5+1) * -1 * atan( 1 / (  0 + 2^5 ) )   n =  5   d_n = -0-1i 
assign v[4'b1110] [06] = 22'h 3FFE00;  // -1.9998372634210344 = 2^(6+1) * -1 * atan( 1 / (  0 + 2^6 ) )   n =  6   d_n = -0-1i 
assign v[4'b1110] [07] = 22'h 3FFE00;  // -1.9999593113858845 = 2^(7+1) * -1 * atan( 1 / (  0 + 2^7 ) )   n =  7   d_n = -0-1i 
assign v[4'b1110] [08] = 22'h 3FFE00;  // -1.9999898275670895 = 2^(8+1) * -1 * atan( 1 / (  0 + 2^8 ) )   n =  8   d_n = -0-1i 
assign v[4'b1110] [09] = 22'h 3FFE00;  // -1.9999974568743104 = 2^(9+1) * -1 * atan( 1 / (  0 + 2^9 ) )   n =  9   d_n = -0-1i 
assign v[4'b1110] [10] = 22'h 3FFE00;  // -1.9999993642174863 = 2^(10+1) * -1 * atan( 1 / (  0 + 2^10 ) )   n = 10   d_n = -0-1i 
assign v[4'b1110] [11] = 22'h 3FFE00;  // -1.9999998410543034 = 2^(11+1) * -1 * atan( 1 / (  0 + 2^11 ) )   n = 11   d_n = -0-1i 
assign v[4'b1110] [12] = 22'h 3FFE00;  // -1.9999999602635716 = 2^(12+1) * -1 * atan( 1 / (  0 + 2^12 ) )   n = 12   d_n = -0-1i 
assign v[4'b1110] [13] = 22'h 3FFE00;  // -1.9999999900658927 = 2^(13+1) * -1 * atan( 1 / (  0 + 2^13 ) )   n = 13   d_n = -0-1i 
assign v[4'b1110] [14] = 22'h 3FFE00;  // -1.9999999975164731 = 2^(14+1) * -1 * atan( 1 / (  0 + 2^14 ) )   n = 14   d_n = -0-1i 
assign v[4'b1110] [15] = 22'h 3FFE00;  // -1.9999999993791182 = 2^(15+1) * -1 * atan( 1 / (  0 + 2^15 ) )   n = 15   d_n = -0-1i 
assign v[4'b1110] [16] = 22'h 3FFE00;  // -1.9999999998447795 = 2^(16+1) * -1 * atan( 1 / (  0 + 2^16 ) )   n = 16   d_n = -0-1i 
assign v[4'b1110] [17] = 22'h 3FFE00;  // -1.9999999999611948 = 2^(17+1) * -1 * atan( 1 / (  0 + 2^17 ) )   n = 17   d_n = -0-1i 
assign v[4'b1110] [18] = 22'h 3FFE00;  // -1.9999999999902986 = 2^(18+1) * -1 * atan( 1 / (  0 + 2^18 ) )   n = 18   d_n = -0-1i 
assign v[4'b1110] [19] = 22'h 3FFE00;  // -1.9999999999975746 = 2^(19+1) * -1 * atan( 1 / (  0 + 2^19 ) )   n = 19   d_n = -0-1i 
assign v[4'b1110] [20] = 22'h 3FFE00;  // -1.9999999999993936 = 2^(20+1) * -1 * atan( 1 / (  0 + 2^20 ) )   n = 20   d_n = -0-1i 
assign v[4'b1110] [21] = 22'h 3FFE00;  // -1.9999999999998483 = 2^(21+1) * -1 * atan( 1 / (  0 + 2^21 ) )   n = 21   d_n = -0-1i 
assign v[4'b1110] [22] = 22'h 3FFE00;  // -1.9999999999999620 = 2^(22+1) * -1 * atan( 1 / (  0 + 2^22 ) )   n = 22   d_n = -0-1i 
assign v[4'b1110] [23] = 22'h 3FFE00;  // -1.9999999999999905 = 2^(23+1) * -1 * atan( 1 / (  0 + 2^23 ) )   n = 23   d_n = -0-1i 
assign v[4'b1110] [24] = 22'h 3FFE00;  // -1.9999999999999976 = 2^(24+1) * -1 * atan( 1 / (  0 + 2^24 ) )   n = 24   d_n = -0-1i 
assign v[4'b1110] [25] = 22'h 3FFE00;  // -1.9999999999999993 = 2^(25+1) * -1 * atan( 1 / (  0 + 2^25 ) )   n = 25   d_n = -0-1i 
assign v[4'b1110] [26] = 22'h 3FFE00;  // -1.9999999999999998 = 2^(26+1) * -1 * atan( 1 / (  0 + 2^26 ) )   n = 26   d_n = -0-1i 
assign v[4'b1110] [27] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(27+1) * -1 * atan( 1 / (  0 + 2^27 ) )   n = 27   d_n = -0-1i 
assign v[4'b1110] [28] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(28+1) * -1 * atan( 1 / (  0 + 2^28 ) )   n = 28   d_n = -0-1i 
assign v[4'b1110] [29] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(29+1) * -1 * atan( 1 / (  0 + 2^29 ) )   n = 29   d_n = -0-1i 
assign v[4'b1110] [30] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(30+1) * -1 * atan( 1 / (  0 + 2^30 ) )   n = 30   d_n = -0-1i 
assign v[4'b1110] [31] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(31+1) * -1 * atan( 1 / (  0 + 2^31 ) )   n = 31   d_n = -0-1i 
assign v[4'b1110] [32] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(32+1) * -1 * atan( 1 / (  0 + 2^32 ) )   n = 32   d_n = -0-1i 
assign v[4'b1110] [33] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(33+1) * -1 * atan( 1 / (  0 + 2^33 ) )   n = 33   d_n = -0-1i 
assign v[4'b1110] [34] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(34+1) * -1 * atan( 1 / (  0 + 2^34 ) )   n = 34   d_n = -0-1i 
assign v[4'b1110] [35] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(35+1) * -1 * atan( 1 / (  0 + 2^35 ) )   n = 35   d_n = -0-1i 
assign v[4'b1110] [36] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(36+1) * -1 * atan( 1 / (  0 + 2^36 ) )   n = 36   d_n = -0-1i 
assign v[4'b1110] [37] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(37+1) * -1 * atan( 1 / (  0 + 2^37 ) )   n = 37   d_n = -0-1i 
assign v[4'b1110] [38] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(38+1) * -1 * atan( 1 / (  0 + 2^38 ) )   n = 38   d_n = -0-1i 
assign v[4'b1110] [39] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(39+1) * -1 * atan( 1 / (  0 + 2^39 ) )   n = 39   d_n = -0-1i 
assign v[4'b1110] [40] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(40+1) * -1 * atan( 1 / (  0 + 2^40 ) )   n = 40   d_n = -0-1i 
assign v[4'b1110] [41] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(41+1) * -1 * atan( 1 / (  0 + 2^41 ) )   n = 41   d_n = -0-1i 
assign v[4'b1110] [42] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(42+1) * -1 * atan( 1 / (  0 + 2^42 ) )   n = 42   d_n = -0-1i 
assign v[4'b1110] [43] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(43+1) * -1 * atan( 1 / (  0 + 2^43 ) )   n = 43   d_n = -0-1i 
assign v[4'b1110] [44] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(44+1) * -1 * atan( 1 / (  0 + 2^44 ) )   n = 44   d_n = -0-1i 
assign v[4'b1110] [45] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(45+1) * -1 * atan( 1 / (  0 + 2^45 ) )   n = 45   d_n = -0-1i 
assign v[4'b1110] [46] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(46+1) * -1 * atan( 1 / (  0 + 2^46 ) )   n = 46   d_n = -0-1i 
assign v[4'b1110] [47] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(47+1) * -1 * atan( 1 / (  0 + 2^47 ) )   n = 47   d_n = -0-1i 
assign v[4'b1110] [48] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(48+1) * -1 * atan( 1 / (  0 + 2^48 ) )   n = 48   d_n = -0-1i 
assign v[4'b1110] [49] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(49+1) * -1 * atan( 1 / (  0 + 2^49 ) )   n = 49   d_n = -0-1i 
assign v[4'b1110] [50] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(50+1) * -1 * atan( 1 / (  0 + 2^50 ) )   n = 50   d_n = -0-1i 
assign v[4'b1110] [51] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(51+1) * -1 * atan( 1 / (  0 + 2^51 ) )   n = 51   d_n = -0-1i 
assign v[4'b1110] [52] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(52+1) * -1 * atan( 1 / (  0 + 2^52 ) )   n = 52   d_n = -0-1i 
assign v[4'b1110] [53] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(53+1) * -1 * atan( 1 / (  0 + 2^53 ) )   n = 53   d_n = -0-1i 
assign v[4'b1110] [54] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(54+1) * -1 * atan( 1 / (  0 + 2^54 ) )   n = 54   d_n = -0-1i 
assign v[4'b1110] [55] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(55+1) * -1 * atan( 1 / (  0 + 2^55 ) )   n = 55   d_n = -0-1i 
assign v[4'b1110] [56] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(56+1) * -1 * atan( 1 / (  0 + 2^56 ) )   n = 56   d_n = -0-1i 
assign v[4'b1110] [57] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(57+1) * -1 * atan( 1 / (  0 + 2^57 ) )   n = 57   d_n = -0-1i 
assign v[4'b1110] [58] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(58+1) * -1 * atan( 1 / (  0 + 2^58 ) )   n = 58   d_n = -0-1i 
assign v[4'b1110] [59] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(59+1) * -1 * atan( 1 / (  0 + 2^59 ) )   n = 59   d_n = -0-1i 
assign v[4'b1110] [60] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(60+1) * -1 * atan( 1 / (  0 + 2^60 ) )   n = 60   d_n = -0-1i 
assign v[4'b1110] [61] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(61+1) * -1 * atan( 1 / (  0 + 2^61 ) )   n = 61   d_n = -0-1i 
assign v[4'b1110] [62] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(62+1) * -1 * atan( 1 / (  0 + 2^62 ) )   n = 62   d_n = -0-1i 
assign v[4'b1110] [63] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(63+1) * -1 * atan( 1 / (  0 + 2^63 ) )   n = 63   d_n = -0-1i 
assign v[4'b1110] [64] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(64+1) * -1 * atan( 1 / (  0 + 2^64 ) )   n = 64   d_n = -0-1i 
assign v[4'b1111] [01] = 22'h 3FFCDB;  // -3.1415926535897931 = 2^(1+1) * -1 * atan( 1 / ( -1 + 2^1 ) )   n =  1   d_n = -1-1i 
assign v[4'b1111] [02] = 22'h 3FFD6D;  // -2.5740044351731375 = 2^(2+1) * -1 * atan( 1 / ( -1 + 2^2 ) )   n =  2   d_n = -1-1i 
assign v[4'b1111] [03] = 22'h 3FFDBA;  // -2.2703528736666230 = 2^(3+1) * -1 * atan( 1 / ( -1 + 2^3 ) )   n =  3   d_n = -1-1i 
assign v[4'b1111] [04] = 22'h 3FFDDE;  // -2.1301812408263618 = 2^(4+1) * -1 * atan( 1 / ( -1 + 2^4 ) )   n =  4   d_n = -1-1i 
assign v[4'b1111] [05] = 22'h 3FFDEF;  // -2.0638004758562509 = 2^(5+1) * -1 * atan( 1 / ( -1 + 2^5 ) )   n =  5   d_n = -1-1i 
assign v[4'b1111] [06] = 22'h 3FFDF7;  // -2.0315754229491265 = 2^(6+1) * -1 * atan( 1 / ( -1 + 2^6 ) )   n =  6   d_n = -1-1i 
assign v[4'b1111] [07] = 22'h 3FFDFB;  // -2.0157063741697390 = 2^(7+1) * -1 * atan( 1 / ( -1 + 2^7 ) )   n =  7   d_n = -1-1i 
assign v[4'b1111] [08] = 22'h 3FFDFD;  // -2.0078328446771208 = 2^(8+1) * -1 * atan( 1 / ( -1 + 2^8 ) )   n =  8   d_n = -1-1i 
assign v[4'b1111] [09] = 22'h 3FFDFE;  // -2.0039113362396619 = 2^(9+1) * -1 * atan( 1 / ( -1 + 2^9 ) )   n =  9   d_n = -1-1i 
assign v[4'b1111] [10] = 22'h 3FFDFF;  // -2.0019543965642979 = 2^(10+1) * -1 * atan( 1 / ( -1 + 2^10 ) )   n = 10   d_n = -1-1i 
assign v[4'b1111] [11] = 22'h 3FFDFF;  // -2.0009768803913479 = 2^(11+1) * -1 * atan( 1 / ( -1 + 2^11 ) )   n = 11   d_n = -1-1i 
assign v[4'b1111] [12] = 22'h 3FFDFF;  // -2.0004883607228541 = 2^(12+1) * -1 * atan( 1 / ( -1 + 2^12 ) )   n = 12   d_n = -1-1i 
assign v[4'b1111] [13] = 22'h 3FFDFF;  // -2.0002441604932146 = 2^(13+1) * -1 * atan( 1 / ( -1 + 2^13 ) )   n = 13   d_n = -1-1i 
assign v[4'b1111] [14] = 22'h 3FFDFF;  // -2.0001220752795539 = 2^(14+1) * -1 * atan( 1 / ( -1 + 2^14 ) )   n = 14   d_n = -1-1i 
assign v[4'b1111] [15] = 22'h 3FFDFF;  // -2.0000610363980136 = 2^(15+1) * -1 * atan( 1 / ( -1 + 2^15 ) )   n = 15   d_n = -1-1i 
assign v[4'b1111] [16] = 22'h 3FFDFF;  // -2.0000305178885660 = 2^(16+1) * -1 * atan( 1 / ( -1 + 2^16 ) )   n = 16   d_n = -1-1i 
assign v[4'b1111] [17] = 22'h 3FFDFF;  // -2.0000152588666729 = 2^(17+1) * -1 * atan( 1 / ( -1 + 2^17 ) )   n = 17   d_n = -1-1i 
assign v[4'b1111] [18] = 22'h 3FFDFF;  // -2.0000076294139340 = 2^(18+1) * -1 * atan( 1 / ( -1 + 2^18 ) )   n = 18   d_n = -1-1i 
assign v[4'b1111] [19] = 22'h 3FFDFF;  // -2.0000038147021164 = 2^(19+1) * -1 * atan( 1 / ( -1 + 2^19 ) )   n = 19   d_n = -1-1i 
assign v[4'b1111] [20] = 22'h 3FFDFF;  // -2.0000019073498456 = 2^(20+1) * -1 * atan( 1 / ( -1 + 2^20 ) )   n = 20   d_n = -1-1i 
assign v[4'b1111] [21] = 22'h 3FFDFF;  // -2.0000009536746197 = 2^(21+1) * -1 * atan( 1 / ( -1 + 2^21 ) )   n = 21   d_n = -1-1i 
assign v[4'b1111] [22] = 22'h 3FFDFF;  // -2.0000004768372341 = 2^(22+1) * -1 * atan( 1 / ( -1 + 2^22 ) )   n = 22   d_n = -1-1i 
assign v[4'b1111] [23] = 22'h 3FFDFF;  // -2.0000002384185982 = 2^(23+1) * -1 * atan( 1 / ( -1 + 2^23 ) )   n = 23   d_n = -1-1i 
assign v[4'b1111] [24] = 22'h 3FFDFF;  // -2.0000001192092944 = 2^(24+1) * -1 * atan( 1 / ( -1 + 2^24 ) )   n = 24   d_n = -1-1i 
assign v[4'b1111] [25] = 22'h 3FFDFF;  // -2.0000000596046461 = 2^(25+1) * -1 * atan( 1 / ( -1 + 2^25 ) )   n = 25   d_n = -1-1i 
assign v[4'b1111] [26] = 22'h 3FFDFF;  // -2.0000000298023228 = 2^(26+1) * -1 * atan( 1 / ( -1 + 2^26 ) )   n = 26   d_n = -1-1i 
assign v[4'b1111] [27] = 22'h 3FFDFF;  // -2.0000000149011612 = 2^(27+1) * -1 * atan( 1 / ( -1 + 2^27 ) )   n = 27   d_n = -1-1i 
assign v[4'b1111] [28] = 22'h 3FFDFF;  // -2.0000000074505806 = 2^(28+1) * -1 * atan( 1 / ( -1 + 2^28 ) )   n = 28   d_n = -1-1i 
assign v[4'b1111] [29] = 22'h 3FFDFF;  // -2.0000000037252903 = 2^(29+1) * -1 * atan( 1 / ( -1 + 2^29 ) )   n = 29   d_n = -1-1i 
assign v[4'b1111] [30] = 22'h 3FFDFF;  // -2.0000000018626451 = 2^(30+1) * -1 * atan( 1 / ( -1 + 2^30 ) )   n = 30   d_n = -1-1i 
assign v[4'b1111] [31] = 22'h 3FFDFF;  // -2.0000000009313226 = 2^(31+1) * -1 * atan( 1 / ( -1 + 2^31 ) )   n = 31   d_n = -1-1i 
assign v[4'b1111] [32] = 22'h 3FFDFF;  // -2.0000000004656613 = 2^(32+1) * -1 * atan( 1 / ( -1 + 2^32 ) )   n = 32   d_n = -1-1i 
assign v[4'b1111] [33] = 22'h 3FFDFF;  // -2.0000000002328306 = 2^(33+1) * -1 * atan( 1 / ( -1 + 2^33 ) )   n = 33   d_n = -1-1i 
assign v[4'b1111] [34] = 22'h 3FFDFF;  // -2.0000000001164153 = 2^(34+1) * -1 * atan( 1 / ( -1 + 2^34 ) )   n = 34   d_n = -1-1i 
assign v[4'b1111] [35] = 22'h 3FFDFF;  // -2.0000000000582077 = 2^(35+1) * -1 * atan( 1 / ( -1 + 2^35 ) )   n = 35   d_n = -1-1i 
assign v[4'b1111] [36] = 22'h 3FFDFF;  // -2.0000000000291038 = 2^(36+1) * -1 * atan( 1 / ( -1 + 2^36 ) )   n = 36   d_n = -1-1i 
assign v[4'b1111] [37] = 22'h 3FFDFF;  // -2.0000000000145519 = 2^(37+1) * -1 * atan( 1 / ( -1 + 2^37 ) )   n = 37   d_n = -1-1i 
assign v[4'b1111] [38] = 22'h 3FFDFF;  // -2.0000000000072760 = 2^(38+1) * -1 * atan( 1 / ( -1 + 2^38 ) )   n = 38   d_n = -1-1i 
assign v[4'b1111] [39] = 22'h 3FFDFF;  // -2.0000000000036380 = 2^(39+1) * -1 * atan( 1 / ( -1 + 2^39 ) )   n = 39   d_n = -1-1i 
assign v[4'b1111] [40] = 22'h 3FFDFF;  // -2.0000000000018190 = 2^(40+1) * -1 * atan( 1 / ( -1 + 2^40 ) )   n = 40   d_n = -1-1i 
assign v[4'b1111] [41] = 22'h 3FFE00;  // -2.0000000000009095 = 2^(41+1) * -1 * atan( 1 / ( -1 + 2^41 ) )   n = 41   d_n = -1-1i 
assign v[4'b1111] [42] = 22'h 3FFE00;  // -2.0000000000004547 = 2^(42+1) * -1 * atan( 1 / ( -1 + 2^42 ) )   n = 42   d_n = -1-1i 
assign v[4'b1111] [43] = 22'h 3FFE00;  // -2.0000000000002274 = 2^(43+1) * -1 * atan( 1 / ( -1 + 2^43 ) )   n = 43   d_n = -1-1i 
assign v[4'b1111] [44] = 22'h 3FFE00;  // -2.0000000000001137 = 2^(44+1) * -1 * atan( 1 / ( -1 + 2^44 ) )   n = 44   d_n = -1-1i 
assign v[4'b1111] [45] = 22'h 3FFE00;  // -2.0000000000000568 = 2^(45+1) * -1 * atan( 1 / ( -1 + 2^45 ) )   n = 45   d_n = -1-1i 
assign v[4'b1111] [46] = 22'h 3FFE00;  // -2.0000000000000284 = 2^(46+1) * -1 * atan( 1 / ( -1 + 2^46 ) )   n = 46   d_n = -1-1i 
assign v[4'b1111] [47] = 22'h 3FFE00;  // -2.0000000000000142 = 2^(47+1) * -1 * atan( 1 / ( -1 + 2^47 ) )   n = 47   d_n = -1-1i 
assign v[4'b1111] [48] = 22'h 3FFE00;  // -2.0000000000000071 = 2^(48+1) * -1 * atan( 1 / ( -1 + 2^48 ) )   n = 48   d_n = -1-1i 
assign v[4'b1111] [49] = 22'h 3FFE00;  // -2.0000000000000036 = 2^(49+1) * -1 * atan( 1 / ( -1 + 2^49 ) )   n = 49   d_n = -1-1i 
assign v[4'b1111] [50] = 22'h 3FFE00;  // -2.0000000000000018 = 2^(50+1) * -1 * atan( 1 / ( -1 + 2^50 ) )   n = 50   d_n = -1-1i 
assign v[4'b1111] [51] = 22'h 3FFE00;  // -2.0000000000000009 = 2^(51+1) * -1 * atan( 1 / ( -1 + 2^51 ) )   n = 51   d_n = -1-1i 
assign v[4'b1111] [52] = 22'h 3FFE00;  // -2.0000000000000004 = 2^(52+1) * -1 * atan( 1 / ( -1 + 2^52 ) )   n = 52   d_n = -1-1i 
assign v[4'b1111] [53] = 22'h 3FFE00;  // -2.0000000000000004 = 2^(53+1) * -1 * atan( 1 / ( -1 + 2^53 ) )   n = 53   d_n = -1-1i 
assign v[4'b1111] [54] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(54+1) * -1 * atan( 1 / ( -1 + 2^54 ) )   n = 54   d_n = -1-1i 
assign v[4'b1111] [55] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(55+1) * -1 * atan( 1 / ( -1 + 2^55 ) )   n = 55   d_n = -1-1i 
assign v[4'b1111] [56] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(56+1) * -1 * atan( 1 / ( -1 + 2^56 ) )   n = 56   d_n = -1-1i 
assign v[4'b1111] [57] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(57+1) * -1 * atan( 1 / ( -1 + 2^57 ) )   n = 57   d_n = -1-1i 
assign v[4'b1111] [58] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(58+1) * -1 * atan( 1 / ( -1 + 2^58 ) )   n = 58   d_n = -1-1i 
assign v[4'b1111] [59] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(59+1) * -1 * atan( 1 / ( -1 + 2^59 ) )   n = 59   d_n = -1-1i 
assign v[4'b1111] [60] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(60+1) * -1 * atan( 1 / ( -1 + 2^60 ) )   n = 60   d_n = -1-1i 
assign v[4'b1111] [61] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(61+1) * -1 * atan( 1 / ( -1 + 2^61 ) )   n = 61   d_n = -1-1i 
assign v[4'b1111] [62] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(62+1) * -1 * atan( 1 / ( -1 + 2^62 ) )   n = 62   d_n = -1-1i 
assign v[4'b1111] [63] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(63+1) * -1 * atan( 1 / ( -1 + 2^63 ) )   n = 63   d_n = -1-1i 
assign v[4'b1111] [64] = 22'h 3FFE00;  // -2.0000000000000000 = 2^(64+1) * -1 * atan( 1 / ( -1 + 2^64 ) )   n = 64   d_n = -1-1i 
