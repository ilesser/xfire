// -----------------------------------------------------------------------------
//
// -----------------------------------------------------------------------------
// Description:
// ------------
//
// XXXXX FILL IN HERE XXXXX
//
// -----------------------------------------------------------------------------
// File name:
// ----------
//
// xfire_fpucordic.vh
//
// -----------------------------------------------------------------------------
// History:
// --------
//
//    - 2016-03-16 - ilesser - Original version.
//
// -----------------------------------------------------------------------------

// *****************************************************************************
// Definitions
// *****************************************************************************

//XXXXX FILL IN HERE XXXXX
//`define XXXXX YYY

localparam E_SIZE_S  = 8;
localparam F_SIZE_S  = 23;
localparam E_SIZE_D  = 11;
localparam F_SIZE_D  = 52;
// *****************************************************************************

